XlxV64EB    3a30     fe0�/�2��cG�1:X\CX�	���;��7��Hi=�<�7�߮�˽t�01ޡ*��01�6k�_��;A����f�x��"([*�_U�0�߂G�]M�V���3y-���S��"�{�4� �W?8{�"���|0W�Hm�C'-���ج���(Q�����ѵ$Ȉ�}��ɉ6ڪ9?tc&�Y�@�o2 8������e�g���t�]6�V�K���:aje�s:�j~���i۠D�:���O��m�N$��l�.���O`.�Lul��|eM$�/B�O�y5FGk��~ݶ�|��ٯ�݅�z��f���^�^�}�m
)�����5�,4�qX2$��@b����#���8�"�Vi���Tl�Z)���Q���eb[�	�=�)�H�9�����LS����1?%��C}&�w�P]�K.}� i|\(��V��G��O8Nl�6h���R'��9��D��o�[Lق\���F�_�p��|�o�vV�c} �;n�,}�E���2��n�֕��,�F���ޖ���q��?,������w����2)�YfO~�)T�D��U��FF�x%.R�F���(�ߜz���	Y������q���G$4Qf �_)ZIzdb���8�$A��n�#��p(V��{�)���qW�#L�]��{��xB"m"3�R�
s�ۨ%Q$~�6փv�(|���vԱ�/�A�_,[���aK���j�Š�MOv+�i#�Ac��,wpvF<�1�s	�g�µl��z�I��@��(M&����H:zB�=��C�[����)����+�3Z�s�DEc+���o1a����P��b�GkWbVI9�T"0�L*�o	jHk
K��>�^������s��E2L�q+D6��l:УH<������V@����`ھ8, �|��KV|T�֝�E���Eg_���(h�����Ɏ�<��ޠ��$N����Z�@��@���^�2�',���6�����c	WU���F�g�V�r �1[��d>+KP��qϬ��J��mԉwF������:5�D�vX��-T�2���Y�``PV��I�P|��@.WNq>�G3a�ը�H�Us�h�y�i��=܀���W�ڵ��K@�hN#�c�΀�1� ��M��pK�����EW)��d�)��[GwdD��'J�nR&��y5��skH3�8����� ��im����,���VB�6��sRǕ�<P�����%2�p�<���^x� 蹣���۩��:��%�0x��9��~�8(����Қ �+����lN�hɵmC#���H��	SI���^��7�3��w�TІﻑ[&.���F���g����دy�C*ȹӅ�ص�XK�b�Sc�}eu�:T!զ������1�M?r�+L�5QtN����-ﴓW|Ũ �J����Qr���a��$�4�#��8}�yLQ�	�0Q��U�J��"�9�������f�?^�>�ֻ�6��+���8�/��ȅ���7@/�$?�|�������:�[�u<���G���+��q�_�`�aF�O_-.a�o����
��~���]���2��x#8$�O���X�[IF���T���@�yݏ�)k��
R6+ �Ѵ���!̄��D;3�I�U�߀���?�^�s����y/��c���G�x�n����,6T�jwJ59n�%F+נ�O\���G������n��@�X�ĺ�=�;%P��F?��̰H�D�v��I.��VhL7KkLL�Y)f&ma.E�}��͆uRK����o���n�
�>:��):�l4�G�����#h�3����C�{���ǁV��V"|���O�o��W_�>mjh-��;55�ϐ��0�'�r͉z�v�}_��@2YW�� �KL��R	nv��P*7;� U!�x���jY]_\���g-QxRÍxK��A��WCG�B?��������#�)1�C���0��B?��A�)Dث�S�k�������g8�f�����PJ��*e�㋷���~�����vy��\@'��m�H�ܭAY��Pp�I�����p6}NI`�
*u�&@^�3�Q���T:~��eLQjj�k��c�mW�#�m���2�#�P�s8[��j����dP����Ӭ!�g7y�l�״H�(�N'x���l�������8�<�񌓿��O��9e�g�f��wg���Q�TԨmt�
��RHY}-�:�0�*����X���BqW��S]�����UDe͑�׫XD�?�r�E^4��i��Il�0���o%a�^�@1#f>��D��'Y2����?��jD����i>σP�w����@��*g�?KOw�NN�x���ܴ�G���
M
�p����+��Ş]h�_��c�D���1f���� �#�Uk�
m�{U:%�-d��tC�Pq�CR�.��Mp� �W�=�SM(͡��<�"���H$��g��Eãy6��LΎX#������On�Q�.P
�H�O��r��fK��gN��;�/9�6?�݋�T�o�J�ʵ�c���<�4$2���qc�,���'*�&Ƣ�<�)�5Y:H8�d��� &�z�k�g#�
,�6NO~6�l9*���*>x�w�+34��x�����r,*�ڜ.n]2P?7ه���!��!͞!oV0}����ZY�à�ǉg0]�_�1Yz�s@C���N�/��?o�)�q�9T���V�Az�]<�����<��S~f����8N���ap��De{V��<	�{Ҋ�����>�k&���ݏM~ r�W�S�1r�у��mx<��� N?A���'G�Z�1�t��X�&lہ~�j�p?��,�6=u����G�j�u0TY��L�}+��)��s�X�����[�x��|0��2�;�u���S�Ȫ�S:F{�dJX���=x�����k�3]��O=9���D)&�@�:����L@��ld�L7�\<kh��C�Ԟô���:dk�����f'=0V�����61��t���l*����O�+�/[r�2�'o&�\&��S3�G�)_��Z�E�+�������"u�x2	{r�!�I��We�'4 �'�J��?>���6�S�ݾ���O�6�Ѹ}Ya����-2�� �@{7�1���?`���"{�Jn[(y�a� I�y@��h��D�'�U^����o��h\E!��>�Rb�M���_TG@.߬^/)��P:���
S	�)O�Nd�n����T�]���+1싧�J8S뻌f���Z/�O����F����W
(��t��uV�dz�*�;�'��S�a�(��~�2���Ra-�,6L��#�bI�H��� ά�k��7#+'oNN���,�ⵣ��
�� �3�4��i�W�����#<����k`��8��T��f�ёa��^������?����m�������q�0#�QX%�hZ�.gR�d�Ģ���G����w���(G~F� �m^�(I�oK���8�@�������O9U�]�o6wzȦ�le�ܺ�b�����{�"m~��s�[>�ۤ�L2��g�?�ι㛿ɪY�0�	�)�<�uP�*$�)k��$�xS�w�񨻐]�(Z�w�w�|��L*a�^���0c`'�5[�}�)�������4N��e�%���:��.�U��޸�C=�_k�� K����-R� ��7�[tGG������7�X\����Dg|Ԗ�\#�DB��Q
U�� ����2�Qa����x�����Ӷ�N�KF�@�P-r�۩#�5bN��`K���P�Y���2=�<Vܥ�j�5b�k]��rs���#������s&���p�$�ˤ���].��׆�r�9�,�Ȝ��0y���޷�.�#����h>�?p2�nY:&���\�!B��GM�Ӌ��"T�pr)�)Н�LRÐG��8�����I���x�ͧ*�/ �m�c�ɟ������F1��'Ap����7�j���zF��4�����Ķ��N�wa��