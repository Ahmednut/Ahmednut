XlxV64EB    28b7     c00�ٖ��p�����߳ \:fUBazH@��oI%�y�x?�r��]އ5I�¬�����LI������Ld_ ���F��>_Q� ���x��fΨH �2&HM�X�`���-�JNd�-��s	�Y�������Ef&&8Ce&$p���p�^-��ۅ�*X�@Ӹ�AqAYߗ�ǘ��嬪���1�
��1��i��VQ�ǉ�v��XF?0o�Z�}�)��-�&�����/�m<o�6ke��l��Nr�ľ\u{wP���?����W!zy��|!'Z�p����ӲO[��K�̈l4?��U��+>�H�P��-N�x@n��x�?�J�V\O=~�NJ֜'H*�=d0�Ps3`��rR!g�R[.sQ9���r�u
cU�X�RJ�*ҷ�y���`��hJ�Ys)m��H�[�� }E�!�o���x�ժ@<�elO�������+ݵ9+�y�rP��6s����\Mc���/�L>�+�^@� ��;<�k��Ϡ�&k f����w�z��F�f�DY�MWe-�S��4mPYfw�/�8B�!�ˈïI�j֢h)��� ��.�2��d�,�IJ�G�K���{�t�6y*�����]�����(m�8|/�z�]~2=��:�R�Q�����mg) -��9΂�pT��� �V��<�K��Q�n[^b�[Z14y
#���"�����h�#n}O�ܱ�&� ��mA�ʝ�DG��%�:�,����H2�"l��K@+��J�oZ}ٌ�����$C��dn�����ܺ/�u�O纻��Ub��5�~�)��&'���oP47L�_@�إW�D2MPb���g�5PMt>2Z�M �h�{�A,���___�3ً0C`�u����z?�L�X:��������P�$�#�Y.	c�f�l�bx�~��2�Wƽ0�S�A�2��H����e�;�ĠE+����.:
�������U��P�߱sm}�Bĵ�~�*�'��2�⿞�ե��o�igě�cI��-ָEN�c�5V������X�=;	��S>Ȅ�b���z��?�2P][C#�����a��{�Q>t�~}�8���0�ʁ�Q�`�XD" ���]>�-M��MQҭ�~ܫ�2��\t��N��Hv@N���m�(�
?6��T0Bwܺ�N���e�#P�:�s8�`��]11���E_
��8�p�����"A����|�r�#�&��� i|��[�	�_�=S8�w�{�j� o�v�\)���E���Bo�\����!Tȴ�jF�Ȥ�fb��o��P���\G�G���_@�sLh�h��=H�������`� �?� T��:k'��(���ٴ�ԥG=&��zs�a���>!0�&���/?�$9���A�"�U90�N�ꖒ=��y�)A?6y"ǀ5����"�ix�	3<
�4X��>��ѸF���
��L`>i��Fj�`�^K���Ʋ��?~�0�-��Գ�*P�{b��yZ ZF�.�J�^uI%��z���'I؁Y}�_��)�VMܜl]�>���h�I�	Mf%⸗ �N�Q������ƕ��ґ�9��w�����0v��$�bb�'�ڪ��c�G-$��
���o�\���ìHc���y�6G����e����a��=Q�y���k0��P��/��>8�dw,�;�(8��Z2�=(N��˽�N(�&��>(R���&2�A(ٰ.f��	���4��(?��z�*� z���e���3R���� �,�	�2��`�j�� E�:��V�<�����vq���d9J���~,鞜�q���d�h.p�p����B��D3e��8���+�����VMz����~�+��=��k~��M��B݄[j�:���	�)�1�=Ŗ�Yź��~{�w%�lZ2��.�8yT�������8��ej}�ʽ���*�s�U<0�D����&��;I-�[oS�����:R�#�`p�O�
>�	� I�45�Ε�
���6i�Tk�y5$��k��/ܱ�����	i^�����-q�W�d�ᕤ/!¢~���H�B�/���ѝt��q����C����#7U�
�����V��Z�����r_�^�t9ʙR�DD�?������'�#��F?�rJz�b��LC1X�9��s�R(��u1���l���h�1h�F8��'@e����K5�Uf�"J]�rLiU=􉏥MT��^�d8D�Y�{��H�\��Rj�Sp��:L�����$Q�J.9���滽|\�G*$���?���}0P|��2���Lv���Ű¶��}�]lo]�k��ne��cKH�C؏5���uq�5����>P{9�@���Iq�Fc.��̡���r�m+��X��w�"YB��ǯ���vi�[~H0Yo$���Ʃ���%�YP*����/~P�2�5���y>%*7�oGm,�0H��54j�#��3��1!\�DۥF���]��Ƌ,��F �':��@B`�2�B={Dc��@a��
��Y΂�a�`E5MD�� %ա�}l��p#�cjv[��`�P�]���J'������"q�)�2ĺ䓐���4���&9���}aHpj�fTK ���2n�χRA�٘�����&`�c$�ťXM~���>p�Ō�d������z�nJǡ��F�g�c����裏u"�wp�-#~�f6�I`}'0��X��,�08��+>�aIf���|�L�L�_Tt��QӇRuc�
�ɘ#��-sZ>�F�s]��EuĬ���"���c�&i믰�e���0B�?*�	�who�5�[�5�}$�jhL#��F������6VI˯�g4�Ic�S�g'2�&�'�ǚ�%��}�"����L@����~}�N b��4��k�0"A��=C
y�����b8&�C���JL�}L���0���җ��d��"2����R�D�I=������!�E�=�D$Q_7a�\�,����;��^�N���8�S[M������q���y9�-�u�3�w�L�/�����]V��D6�n��(�m�m�p��c��4�]S;����, �:#K��