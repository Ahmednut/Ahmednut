XlxV64EB    295b     c00.VL~~V�s�%rGA@S)���1ɕ���q��o�G�g$۩����t9�*W�u\b	
K���F񆳘E��]���.�bZ	��nLÉ��+����V�c���C���ڐ�u:Gn�x�5_�Sss�.\����:f\�?�&��;:��ӆ��|��v+�����1'�F����
�>�u���{0�|
�g;X)���aM��+\��(���b0O�ګ�}k�9��UI����=�枋�k��>���YRD����f�!b/=����ZlY���{�|] ���Z�#Ba���^Cf���Y�����rϬ�sF���4y"����=.����C���ςk*ػ�%�G�-�N��я�@�'@�15��V5{���y�-J ZMn��߯S;,�W��r�&�B�A��� 1�:Sj>6��^�����CބPMQ���8ƪ�7$���f�;e'.3kR�ؐ��H����sy�D����\B[`�f?؁#�D"W��`��"�4
�A��8ҧ]���u�#�ks�Ұ��7��o��5��JEj��?��l��X�U�[L}�&� Q�O��jp>�se��d�#2Kx�f��F��8�D$")�W�	�/�i��e��E�k�l�,H<�p�ۮ�xK\������-3&7��#�*�e��_h�D��v�(�J�u�c`sr��,�5Bsg��7��ڲ��)�P������cc�tH�ynM�
�Q�At�����H2�z`E�I;�q��8\%��N�+{�ހќ��.�yH/�n��Ю��:rh"�0������O�0T�K$�+)����J>�@��G���?O��xx⥗�,����6�`[�_�Z:>�Gb�Η��}V8AD`���H�,��A39��v��?Q���
��Qu�)	@r a�ӊ!6�#��b�[�mM���J:ʨ}S�H�U�qS�m:��I�l��!��߁�d4�a�E�������P���A�{&]��Zf?㵽�PҬ|N����p(�A���ΈS�������ޖ��O����{*���ҿ��x���iȻ۲� ��=8�����iQa܉֝6J�X��Q�l O&�UNw��\�=u�;�b�jW�c"?�B+}�)�(�uEG��h-�k�������RD��]�4]i�ZC�SXx#TeOdG�� ә��`�nw[p��c��2&���~�i��ξ���6��#� ���֥/	nM��c`�:o���j��j:i5V��9�S�17�@�O9��0ܴ���p�b�Q滕bm�Q��P|�/,��*�
=a��	�}�
�u�'6��dY���8����!sxմ�Ã��p�H����~��+��? �ƥ�ſ�@�Ҍ�<�@���TO�<(
����Y�}]t�<�eo��H���(�u��ژ���>�M�!3��S��������������Ρ����s������Pf5�{ѥ���G��6�@o�烼?���6��W��Dw���X�)R��2�q�"ER���.�L���T�ގ#��R�4��m����c8�:�{��儮��5�����'���%~�g�~XI*Op��ER�J9��\���o���4S�� �,~/e�Q1���%�4��k�rS� ���.����7�U:�n�>��q�D8d8[�	�
��]��8�D�A�2V�����\�y�}�dx�'��eV/��BY;�\2�.�������J&Sx�Dq��=��.�5��4�q>�J�� � �a�w���*X	��x*�KLRv��ҕ:�eӷ�K@N:?������&�v�R����m�����V��p���`�(��i��p�oܔ�]�٥J�'3оk7���Vѹ�t_� $��Q�%(tt��-=$Z_徝�,�G�U�骝7B���o�?���>��!�C$H�D��ndND�d�Y�Ve���y� #達�g��skzyR��[�~<-l7
�&}��aW$����\�w;��&f��v7�J��b�᳉T��L�~+�V�ъ}��WGm�������R�Niж�&n�)���P'(�|�K4�Ū��1��6^�Kk��PC\�o������ֆg�#j��.ҷL�����f[�-���'��������7q�٩Y�Q��u��f���_�����[�����?X��7�w�~W�� �G��l��{�;ش��]b�4m{$9%�_�\)/@�'
D�7�9�`_*i�h~��>]�w(��<�gz�a�Y	-���޲`Yi�4"�=���TO�>N���,���z<��%�5��������/8-#�5��+�EB���t"�.>�G���&�[�c��i�ƅk�Lx�DA�8�4i٤��]�`�W�DX��Z|�Aa)��C3b3�$��m
����?�3Ȯו�)x�%�����f�c�\��#X!�萧ߓ0�w)�K�k�6�f�j����£���K������WKuE���b7�u���x1D+1&.��*����W@��� ��/���&�e�-�v/8����z|o����L�)�.�7�aa����/o��N�V�P7���99�}>z�K/���GG�<3ST0;�y+�Kc�~i0�	(5���P���j4�wտ�������0����z�S�)۠7,�����F���u#b��i���/���d׎S�c|�C0����af+�>lKKr�V^"�~���7I�Y�`"|E/��Js�U�l�(VF�<��,���.�ʹ�!��f�M�}��+�W��BZ
�@�F�i� ��!�'���b��M�����,t�ԛ�� VN�/N�M+�j�JMS	&>�����0P��Q�z��x�����D�o��Q�ԅ"�wߜ��^J�-�MB���w�p��}����Ȭ�]�K
��=�f�gW66x]|kDS��?R�ÿ�?[2ſ7�UV�+��)��>��
�C���cܨo�`��q�;
�F�F�ɵJ����#o���݀�I;EH3R���:�J�r�ñ�(>O2%��