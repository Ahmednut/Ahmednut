XlxV64EB    57dd    1340qɓ_0���_AC�p�w>�6f|�P�H��!_$sY*�w�Ή�:��Y�����,��=�K�23�q�������,쥦4�4�q	�� ���8���SO<Sc>�C�G8!	���̙\_t��v8��-)���4(�.���A�YK�:^��_�P�=��)�v�&��M�xګuy��lk�"�-�1*�����J���r��q�φ�.y$j���NE��E~Ǘ��� �� J�2J�%���j���&�ڱ LXH�9!��O�O��#K�^����8e�q~y���5yN����-?P��{4Z�v��&�hl��Ű��Ӭ��"�"9���fQN46�po��F+�2?gA�ԒX��|��1Q\XT�!���#m]׊�u_gI�Mu�>�wFԀC�o̽�ϬDE6]��`���}�W��m�{���vV'�D��b�8�s J8�_16\U�f�TO�T�g���C������sk��=N��w�}���rb��p��W�;�l��hH{N�{��Wk=��֘��n{ԒR;����}LV2t��3v�TJp~�q�p�'���;�@���K���I����֢K�s���Ga�=NX��g����h�'��)FC0�)���'#�;��EGU�6|͢yD&����	�_�=&<*n�~��c��˳���Ȁ����gy�'o����4�o� 4����G��	5%���[�+�Rv>7�8dX7A�Z���v<6�?E�4�_�?e9��l�ꜚEe��B�~ɢ����)q���tD�^L�%w�#l=e��Jn��ʞS2aQ��~���_�acx��� �p���;[��ĭ��Mu &]��AN�cz�{16�M�NR�S����	ڣ�����U��R��R���Y�P�7�3�dz��&(c��&�բ�"�?����#�~�<�c��+�b��Qul�r����:�.c�*����k��O|j8KͰu�q\��|2C�3�\Ob������.b���*Le��<��˙�nT7S8���|�K��V{X�N`>BB}/A���0ǎ7{b��i.�k+R]�)=7�I�[�\�|��t�I��%q�Z�HQ���(<���M4L�Z��~:���X� �;"��{�`���%�n��o�����g���<�*�W��k�,)\��V��\.��-3w���;>P��"ὖ2�0R䱷:�B���įB.D3�-}do�+��P	u��F[\xG���$��L�Ap�a���T^ێ���"7���k��m$a��.���ݬ�w�鹨�������ԯ�nu NGsaZ�>2����k?�����H�Z��E"�y�&����Qz���"%��=��tйb���3���5nty�g<{���oqr�d�[����� ;���@�kZR�ǂt�u������jI-�����_���uv�AC��J!�����:�}ݒ��2g'X�aE�6D�GyC�a.��D~���~W���{USW.�1�A�J2��O.D}�r�<�(���!�FFw���s�>�t�*J��a'%p}��~x��o����˳�P�Ĕ��J�<�H��cQҲ���V�|�x:d��T��5M"�["��NO{+ͺ�6�2���X0����(-�L�sM�w6|��Z�)�R����:�?��������o�UJCU�
���p�;-t��4y�4ЏP*qi5����N���6#��T)�m��R`qV�>���P5?)�l$�s�cMI�Ξ��x��s���&��Z��z��p�v��Eˡ�ӹ��E�ב��7~�Q�m䈯���]遃��v�Gl:��,,���`]�t�mi�J{��S޵��rK�v����W[��v��n�[z�{k�ͯT{�w9p���?^���"����45���VG�����^��ri�VHH�Y�d�� �鮹�n��2>���k_�\ш5i��R5�cB�@3�*~i_d?T�(�o�N�	�
�bO����p,k�-,��"=Z��<M��N&_5z���F/;m0��c�&��L��w�52�Y�N�U�D^V�ڼ1^Z�f*�LNm��D��_�u�K)G�>(�? CM2�2'�t>j`���GIgK��Ƞ~��Q;��*t~�7q�c�֍�k�V�2�y��J4&<�<.y>�Î�N�]W襅�~]�|���b��3��]�+���uR����i��h��7s��/�q��dx/�MJ7Da�Z�gι�%����;���ܣJ������K�D��� u����~�i�U���B�OD ��cɮ�NP�	�͝�"Ѯ��#3�	��[h������y�4�.f+K�w$`f��z�W ]�i��BL�9	C3ӷ�M�֠*9��k�4s���� �/o��k��솣��`���`f���z�~���\�\�{	����Zp��
]x�g 	�V`����;��|�%��{/��'.��GB�V�c�¦by�d�(��z-��� �),ה�
��VP=���Cb�]-/�C/�S&}S�C��B��L ѣ)���?RN�"�'�K��h1�D��	N.��8}��2�r�q���y}��ۜ��>ɮW�Jd��K����k/�����e1�*��_���7Aj$؀��w���,��ʨb�z��V wB�p��$B1�iM�-�-ܭ��m'maLd�Ml����%��[���C��n�6��<�M��tDC����=\��C���W-�cG�]�|+�o|�f	�$Q\�փ]��8�6�՛��j�S�zl���W��S}�g�Q?u����e�(b��:�Y�V"����W�+:�!�_J��8!0��Цi����-�_��WE��U�ӹ���W�`��R�Ԭ�ͣ5��<�g��a��n�1Z�0K*, �6�n��&�8�Ԝ�% jV1�#������� ��(����o�I�jw�D�a�Q���喷����`1}[aI���q>�ԯ���k#�3�n���̘��]rX��۳��48���i�|y�+ǎ,�􉔏`Fڱ\���Q����{y�+�(�X���{M�l�d��,0?lD�� ��S=��%{K�����D�hz�-���	2�����[�R=�E�x��ό+Xki��-��)�M6�k�S����,8���4X�g�Oګn��.iOe[P�*��nD��e�����Rң�����lx��;��kI�Qp�,���a(��x�t�<���y��o(h����e�M�e7�qm��2j��Z:Q��œ����>V�K:N�#H�z����s�����'�u���C׈��3�]~�����QQ�	���4��;�<\�z���%S�x�[rƴ6-���?'S�=�:���n�<'"Ήzv�ڢsZ��U��Z��4�5��.���e#8��I�P�o�qu��/i�օ�ƎQ���[�%�U��t��_�>�/�S�����k��0r�8i_��o�%��N�%.���}�����kxF�R7�)$�.��s:U�(��"�K#>��Y��S��+Xp���]�ՅC�,��9�r�ƨ��#�3�f�d���v�G�	n}�*׿��{^�������AE��n���*i�5D  ���C��He�ח��T������,���K��l)����Q*Lzy�:��&=p- �S�¼����-<8b7���N�=�O_���v�#^Ps��xm�m��|'y�s�F�q 7��j��ďĨ\E���m�]( <�k-�Q)�B�cv�L�md������g�_�*���9��f�!�Z�ڄ�v"A�s����*H��0-QcLe�^t�r|�4��J.W+	��MPfTJnۡ��Od�v,S0�V5Pi��� 3!��V`�t��F�Ȟ�T��yo6�d��L=^�yU�.��A��z-yqdtd[&�ŗ��5��+�:�j:y���Q�
H#�����o��K�ݬ9���w隷��!�Թ3���G'��_��?������n�^]����0\���dӇ ���(X�ije������!3�U`�4=�k���4|a�m��l����2SX�Si*^O[��?ᄱ�l����������0#i���Y�qB:�'�s��^�=���8*�&%!�9K���.���=x��#��օ�s��޸B�_��C���d��Z�="T*E;䠍/��ׁ��0t��g�~\�:� ���Sx��\���N�l�Ӕ��δG�LD<�Χm��Y*X�(|���B}�8�?h���اܔ�ed�}�T�@K��ZK}Hʩ%կ�W����b$��Z*��t��=�?^�_~�gK��G.<�6�����v�Mnr=F˲�YK/ �n� ����4�M�;�C���巟S�����K�gڿ�B��Ŷ�����M��,�C�2}h eafz����Ԅ�� ��<"���tj	��a�V���d��p��m�Z>�0�-x1�u�ÔӮa�XC����J�Ea�S���o�m��s�`��m{ȭ�@�p��@�(��A!��r����;	xs�Jp���YPhW����9�`3m�X�*#�x�����a��������K�S0����t����%}�Էz4Gwx�{��?���w��, ��I���c��<��\E�V����Wc�7�F�S�I)>m�S`��my���[���Y1j�Pӧ����UO�����׋م�A�����#O<�����Fқ�M�P��|||�eG�]?�gep�1�
%v�1d��*�R
�;�KJ�9�q�B�i�wx-�	Yl �LZ�9���?ʜ�M�ypF���WL͝t�:�]sԕ$�����k-�QE�v�ݡA	DAT���[��?�p���I��E��!��6�