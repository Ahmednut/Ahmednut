XlxV64EB    3ba9     f30���yXp��L[�P��^ٌ8gLR����;��٬@�2�s3n�B���حK��^�G9	�R~��WN,_A<1ܷ�;Njs���L'��.�5���#�*�ޭy�
�6�����^9��jB�Z��_�\���nA7�ޡMƨ~n� o'�>A���x������N\"�[O{RF��}ЍM��n�[�h�p�]h�de�1��;<�Vt���w�ڠ��G.�T��H��7
�Wg�k����]2;WW@Z���{a����H�۪�f���j���$o?=�:9@�����e�9�onR$�� Sl�����k�{�m]��� 7-��%�����3\�3F%�|��I֌�ZD��C����%Zw�-,�����8r�x�f�����B�����8wIJ�굒�B�b���J|lc�fj�z�p���uAo����D>�h�s����A7dfh�j�g�u��~'|F��嶤n���8,IV%�V������R�hQ�nļ���&2j8�ᘯ�ca:�e<�߽��@�6J�(���G :�S�E*���+�W��-K��Ѽ��������x]��aeߊc��|��iXSh �t۰AB�5��3�>�U�j���O��zբ�z hE
c��H8�X��.�3��-sv��(�;�$F��
J�t�0�TU�^�nF���,!���N�*Y�c�i��-~�h��k6���_R�sFPpI>P�6;sc�2��ض��e��?[D���H�}�V?�i�|?0�uV�
�h�t9���k<�8�Tz�������;{�����������߮g������P�ݪ"H�Rڏ�Z��U����;�g>�Y�r�5\zN���
�������== �4�Ġ���G
��.�W��]A���C,��D\5���.��e%T�!���8Έ�Q'�ގґB�=�ڭ�BbhM�N�s @ë]maSʋ���淩] dU��.4�R��,h�A�fĴ��{� ���.8����jU ����#� �;����fd�.�P�J��ۂ�_v�����Q[�҉���%�r�Rk}�VK,SNC�`ɓ\�i~�*��5������P��9�(;0�Y ����L.!����+2�R�{������ê������-i{���ڒ|��|1���-&�όN;>�$%��)X�	{�3q�)ֺ\�f�EG}�&��OD�Y���J��SI��n��V�!)�T�`np�Bl&�6�=�MO��a��u���XG�Z�n����e���>�N2�S����lװ�A9�FV���W�]�tK�ZAk�r�%0�J
� +��I$�ێ��ԢL���=�����-�����Ɇ��`�%
y�,j�r����݅=F����M}����@f[�tp���,��
�|�X��tR�:��*��4Cb�%��ɇSd��п��1��@"���f3?-�ű��q
G�� )]G���8$<@CѦ�tθ,��QA��?!
�ڽ��^�	ֿg&��{��(-���mD,q�����dB"��3�]"�5�� �z���jȺ�'��챠�3�U��
	P� $|�� ���Y��aes~+�_���`����Q��:36�-�Ef�S��C�Us���^�w
Ik;|�s�5��_��	5�M5S^�:��uʩ\��N�O�K��~	M�ϳ��y_��ө�bC��y̛*�H
���Q�cꄺ[/���Z_h���F�ĮvV�f�TƆZD͢4Υz�ώ��)�#Qɕ:��r$���HK�k��a�ЗfEk��vB]�
�s&�S[@��,V�q�NɎ2s��r�I�a��*B�a��em��|{�W>u�,X��d`c�b{�.�ۤWh)���n�q���=7���7;Qւ�	�AT�ٷ�g3;�E~n��}� 7N�m�e�L��%��Y#D6h�FP�$&�~�1�n'�!FZ�=�N���q��#{R	�bR�&:M�M=+��x��[E�
�r��^����LU�/�����}�,���J(�f���.�XÄ��`c���7�\���O�������ͱ!��l�Yw��[��V�����9���D.1��n
���;�*�8	�a4��=���C�Xa;j�S<H��v.&�f.�V��:B���g�׀������Ϩ�!���n�6�yqC�CQP��•K����a%����^ft+1)#�����{�]H!�|Q�k�?aX9�_��G��㺱�G�/��qϧ�u	�b��`CdQO]������Wj0��z�]uHE���7�b��k=��oZ�Bo��P�|���l7���.jL�8��C��f��L�V�U�ps�� �<Zh����2���pD�~U�����kLف
"��웕����ԡ#�9�L|EW�qG:0�g���8�v�b֦W�ȭ�ڢ�Ԁ�WKW��H�"0����"�^��q�'�vaҫ��>�4$���sAj�UT��3�LQs{���^�K6 5]��Ý�B{�=(rV���^'��ku�3�����K��w�)�]���, ��P���[�'��˹L����/���m��E���D3��聨���u���T�W�8�t'?mxM1�y�O+*�}&�5���u�l���A�o�W����k�DM4�h�>�-�h.��ï�V?���h�U��ʗ���w�x^�i��ʠ&��J��Ɔ��+/{[:�2�A9�q�-rO�}���\=��������({P��m��4,��z����~��lDK8b�A͘(��r>约�L���A��KD�(��\̀�3������냧�LǕ�P�ڀno^���j�t5�K�=��4�`&��� ��<�o��]1�"M7�pG�dqf�ro���Ϟ��"�i�yU���_}��.S�N]ܬrcr�)�&h�Rby�b�goG�b�qB?(��8~;��n�%�7\O��'s�F�~><�R��%��
kK#��a{Df,�Ѓ,��U*�(Y ��Ϫ)�������B����=�**� �q�޸��N���k(�@(��잿`@ۨ/	��3t,��{�ܮ$_���{D����3OB>����b�S�K�!LNL�Fo��|4{7�@��L�զn���}�H�d�(�,���i������`
*�Wj�`u���tϧT=T� 7QEܼ��tnOpv�;I�ԸA�7�˟��K�7�0��&�0[�Oc�|�Hk_n�I�Uh�??����te�d�YըN��85�߾\n�1�m����$�̀}E�30���qlE��r���/:c���pqT������ �ƥ3��r!\����ʉ;���f��y'X�|�%�%�C<C}�e!N�i z�Q���i�2"wM��:��j�#����IS��m?���;sF�5>Zټ��(P.�*/���?�i�]�jM$��1�f�������2��nׄ�B�8y�1�'-�Q�|����(v�K;��đ��dŜD<���p7Yk���-W<ǐ��
���frg%��'aD����oBi�*��A��R�Op���xI����l��Ly؄�� �ų��S%)���5ԑl��V�Gǰ6$v�"O�õ�'\���Q����]�2]����R�d-�}�� h�3�i�B��~z��%pV�kV�z)�iAւ�	�_;
�ʌ����4#t/H��f�)_���/!�_L�3���P(�Ml�[�����S`�6�W��2��1�u1Ն�������1���c��k�{W�����e����@?�x=�`s�l; :��\C%�X]�Д��^v�p�H&Z`rj��/��k�,M�%���,��uf��45