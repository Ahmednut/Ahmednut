XlxV64EB    7a1a    1a20R�)�<��55ɯ�aJ��
3$���ܟj-��Cؕ�?v�3]\��:��x�ĸ>�9�dyY̷����_���@�R���!n�����e����y�r�L�4	�%�چ���x�=��7�zEO��B���HG�ىN@A��� [��)
��J�� ��wY"L�|��]����6�g����/W70��q&�ga`����	�	Y	9�ӒB�݄�&͢C��΅��K�l����>%�4AK4<�6�����I�R���'R[׌%$��6~�̟p��c�wD�����Ԣ��5��[e�=�Z�i3���ը�X�iӢ�$��N8�ה \6�	3C��6��JW(�`��*!�􎺞�_:m�q���
��樂��'<{�_Ҳ�~����y�j>�Sl�wx4��V�f�
�z]b�F��ި�,��66�Y��o���=����HN�M��;���E@ƀ�G8�+M�^�m��t�G�tN�A�U<�:��5�hW^�n�j"=$�j0; @�B��ˏ�����?#J:f3a(���imC�g����M��W<�kT��M�XItb<�,og#�*8�if��Mp	��n	��4�Dxs���ϙ��th��L�*`�/���I�o�C.!n>/2<Ie��Iқ�q2ͯ~��x$30��œi��{.��ז~:���fN%z_�W�_��Px��h��\��Z���ÈId��l�n\`���U�"�+'+g�O�h�ī�a�@��d�6�T�sakP�J,7s͘�	X��b�7z&�eJg�z�C|s��J�%5�������w|����\�v�,��z���]=:��m[����9U�1%`�W>E���ګ��'��H	j�d��Z���38R��y ǐ�0\����5*�_e�fN�!w��cW(x�.�bcwz����0`ź���=.i�>(7��d0��t8���p6�*�s2+�B�ĕ*�gA��~4�=rq״���8��W�v���M��5Q��9ݬ��XW*=�4�q�@c��C1E����=V���+�'�P1d=Y>l�:�\����Dg�*ƽ@��τcF	l��/�0��kI'X�Z�(���ܻ��m�hN�CZ,��V�57z�Q���5.\�}�^�o�7:A��Q�Kw�G�9>��*�9��9��]^@(�����	��=�@}���l>,5.W4>�U4�H鞘�h�Zja�y2�M3Yj�l`?ޜhxm�jd�ۤ��y�9!3�g�ՠ���R��V���]���4�.��~K�ک�h���\���we��Z���S�z�>K�&�f.��J�u��n%��x�hj�+
ˀW�ͶS�ޚxJG�-�u��Y�y�� Y�U�Id�,jB��p�)�Dp=�!U��0��=ӊ���I�!'W^��ǵf
��g\�8����M���6:��;[�8���e#��Xה��4Qq"K�&I2�Na���]@�m���Eb�)�E�?�fE����5f�`�)].�D�iRӵ���#�a���^Yd/a��b@9��Si	b����b*j@��Q����^�l�u f�f.��4p�8Ν$�$n�DA�Wn����4^��|���6�oe���Z�RZ$�������-XY�*h� [v����Vŉ�\J��̆g���T��ī��)�`�Z��k�{k�1��E��*���Q��bX���+4<�N���6`��wyy�[�ޜ���TU�Z>+6�r�����·<ZEni5���sU����mv��=�� �i0������?�=!���%w~d��K����7꒥A;�82R�m��E@�!��A��
�f�a':���$;��7o�Ι�U��2ݢ���� h���L ��*.?�2ݽD4��
�i�����`���<�q�c$�%��pT�{�B��6r&���U��I�w�v\7D���]��g)��`��e�r�5�)��o��7e���+/}��ɭDu�$���y씿cC��Bۻ���χ\:���"݊c����_Q�����ue�-\��
P7����e��M�oƋ�Z�I����:v�a<�)�O�:�g���.���:�D5���K}����Dt��m]2���&Q��$0$�A�Sk�.2%oI��t�0ɧR��&��	�	w��4��,%�~��ai�L���YM���ҩ�������~��9ݣ��]i$��O.%ŝM���+�	G5f��<�r�~�u[��(?|y��?���@�>
��&�?�Fˮ��A���|�i3��;%���¬\�oU�ٽ�T^J[�X8b�>Bǡ��@l�Z���(�e
���rO�I�����HT�����<�{E֮��*�M�t8w���UB7�Z���އ$���v��e�%���0V`m� 3A�=�&���+a��+�ˉA'���&���#o���R�M�/���8dʟ(-M*zz<�9F�f�U�����FZ���i*�/���:߈�%�����s���hl�\籕�@�c�j$��,�_az5@#��il���3>+[�="�8zDv����	a�\���>��ؓEZɭ85 �^
��j,`WҶ��[A�����o�u�a�U����C�ӮO�xVi#��y��W�j^fV��_��!�f�yk�P+��E�IC�/��	J&R�	=�X�����x�Xk����1vl/���Wg��;��c��X��/�H�DW�l�m�J��n�V�n��ئ]��ۃ��N1�ᠪ��m �<X��9��8�g��p��R����)S|�`�)>S����%�r��X ǉ�7ip��d4�9�s�|a�D�m& ���f��I������N��QzxQ9.��ڻl�w�_�ؔ�]��Ťڈ�_��ȼl���
���aϤ`�.��E˖�9�&<����@`9c(c�*�V�a�?S𱑽�-�*�ّD�tq�u׷��"�'`4�����(�J˒~]�78��c�
I�1u�[�؎�����7Q:�ޞz f=B/#�<���=���!�e.W=l��LS������)�~�����\DM=�,��n�rN����(�SE� Ts���|a�3�p�5���V1�#�|��e�����:H�hC��u��EX3G����5�eih�k�� ��x 2
�m�z�L��%:�W�/��qV=d�2'�ۘ�W֭Yn���V��kc���/��@30��c��p�^���M����R����F�����7��]�i	�P�m�F���s���+'8/fYԉ��!{���t��yyK$M����Ę�>Oñ5y�ۅC�)S�lF[����jX5�ЧYV�G�v��Cr�u=�X�6sxK��.ym�]�&z�x*�ɯ��<"�-S�B�;@1�-.S�;�[����G�����E�y	Q�\{���]���-j�S����Û���rY�DX3qkԒ�5B우e��׵�T��Ê۠}:ֶ���C2[Rg�c*�NX�竂�*�48��3C�Xv3��r��U�nr9���&��|\Uo����PZ�*�7�L�d�<,w` O�\&=n�.'Se��g�!X�JBމX�v�8f���BEj��f�jH'�	kTf ����H�� _�c�.����e��0x��ҳg��!����\�����ڦ�I&�����o���
mU0b���v+��܍+�aaN����EX!?Dvv�B�{&���o��>�� [���;�'��p5l1k�\�����y��lx�c��.h�4%�)r�ƿ�����0�%Q'V�~0"�s>�\j�c�̓!�6|A�2��E�k�V&�<g�D�|���K4��9��Xy �lڡ���(h�Zh�
�G�H����U��k!�aާ� V�/:V�Wu��ҭ��6��W�#}r{���D�0Jj�,����$ē��Ph���eT�5eyҸ�
k��0���)_]�(O�Z������|�G��#�*�w�6�
�}�6ԮE��P�����l�Q��j+J�姱��.g@&j��Zxb��8e��(�^h��F�g<���,)޴&���~Y�F�.eQnzi�mFO+d��7������4j'[�iaK�5.�U 0,���pI�r���}#7���Ήw�ƥ��¤Ei��n�����GXi��Ƕczːyhu�Eg�ho���H'~��|�pi0�N���[s�*��0�6�(�И~�#:��F��6LE0��->��Z !����i�s�(�cPzu���
Lˊ�|�C�kӈ?P$!���Qd�7"��c���y�D�-�A�ֱ2@�o5y2<��V7�2��"�y�C��k��9�8 ���,�"�6�m���`��* ��A�4�q2���U��9ϡ��:z��I�R���;��B��H7Ӱ��e©���J&B� a?���f΋��Gu�(���q���ȁ�A^��l�6}s�=����o��D�ru�C�s�����r0�nWؔ$�~����v��d�d��0�
��w��V!�١��b]T!%%6�XjU>���a��(�������Wj�QA6��q�ȅ_?qǰ/0�
��)���bg�|b7| ��z25,��rCWgù�C��*�W��!X;���rl�H3K:y:b��n8��c.���TK�:�'�v�ג$�B?��H�iph��3��x;����@	�J����E'k�[)?fmG4�s5�>�OL�G�;:�R �g�l��=� ���ř�~�����&/���0߳��,�V�
�����3����m���>�Bwo����x�����}�+��n�!t쌑�t�Kp� �S���6�w�|��76f��2m<�����ʤ�1#nl#2:Ap�'��J�[�:dMf=LC<��,�0�o���{[r��[�Y&��	�t�}�Uu$����dl���ô_���tP��/��J�7)��\��$�\ɍL�I|���E<dbգ{�/{�^��9?B.�H�~+tʤ���Ʌ7��;)THO>�1=���*�]���P�i��Ƽ�ϝSSF���~�8j�-�@��F�D��`�=>��J��s��>�:s�X1�*.H��3����|-���]X���HT���(����gJVo�#�� ��O��i(���~�B{���]{�TE4/K}9��f������N�4�7�U>�}W��<n�a���1�v��@���l=/�}-6}��{Y��4*'�F�@���PB�0��D��5l���$�,uc^W 4ב��^
�Ѕ�Re�{��,�����Z=nM@�%y"`Ft���8��$ț�R*D�N[��J����
~AZ�`�5�d���c��Z	�o°��(�IJ�v���o���o�ؤ'��顯]����*�}��/�lF1+���A6x�X�{_�(]��i��a�~p�ȳ�ݺ��{f��pl��QG(�/�	i6�)\��
����O� �?G��1T�n��v4�>���{wP�9�:�d{�����csu�a.H��k�E�Ndmtgq�VκD �cZ��]�)��?|^��1�H�X�M+�c�x[��8������	*0�����"� }k���w��!IE����v��^�
4x GY+� ���6y��s����e�$���D��K@�@�&��7WJ�p^��n��3�f�C�3�桀�P�0��T=���S�7b�I�e��k��T0���1�VFw�-P�7FP鴴��>�Nk���Q_
���W{�£�	+��л���h�kiA�5�qe�'vO�]��<����K* znS���љp�k�ɀ}�1�Tv\uR1"Le����`3���	^r���Y��LbKh#r��5�YEK@����*R�>�qSա"�jM&1��{\�}k�}�������4J��z����.bí逦��������)�_j�{�.�E^�Y��+D�C����#1�ny!�X�AC6���^<=B���ٞ5.:~��B(�c�_�v�.Ʌ��`�.wՔf�ū�TTp�I
�	���'�"�+���U�vJ=�%L���i6��Axv��� �Fk;���W�`a�J{�U~�N�K"T��4E"b�eC����:0��>8�R�0j�"x�`1������ܜRt}�Z��^J~.v�I�I%eJ���oS~7��1�D��bv+� �T(R�S�@�K�Υ�[��lL�hJ?��ˑ�%h�=ҝX�E[Z�Ӛ��~�U�*ةi����ȷ]r��Z��A3u�eTV���/��ҀZi%?a+�{�f������2+�>r�Ս�'�׫#7�wC9������
��t�m�0�3c[�]�M���P��7P�`��0I�<g�I� �DO��)�[-�ꓚ������_Cq��u���O�G�a(�I���켹�ѫ���/�E�I����!��Q �[����^w U��J�
HFV�e%i:m���|rN��n�)�kم>͍�p�'��;�v|����=�rB�- "��
ܽ����4�y��V�0ޕ�E��V�]������5�Ղ>%hZ�� N��w8�q�lA�N���(ؤӌ7.NF��m;f׬��/��D뛬CoN��`�*���7ݾwB#_	M��@�)�KV�&����