XlxV64EB    fa00    2d40eAH���������*h6�Zt��>�rL�2?]�$�i�}�+;�7�~"R_o' ���q.�T?���}[���k,�����Zw7>��c�лf<lCϽ��o���X�O����3�؟hd��l}Q�(��u������GR��BA塶�wY�:�v3���Ql�B��;u���I^�:Ι+D���g�3��b�ρ]�����,7p�&HE��J F�$ʗC_8A+�i.�c��'�?,���N��6]�P̺��F�V`�e��Trr��;��� �ۃ|��S��绋��=�g�Q�;Ӷ,x3�Ť���w�-�0k���4�1�7Io0~�YS�)�rVt���&��Mo�0s��굵mE�G� y:DS̃�8mÀ�'�`��J��X�;��=�O&n���ڞSk�_j9}���[3ٔ}�n�D��K�5J?8�~�v���;��ػ���r��%��wg�>z����� �{5�8ެ��'!���2�g-'Y)��X*1 k$����u}(��-L�b�1KJ�1p]C��_����6���.(�]��ћ�:wߘg;�9ҝ�J_9l�5|)�)��1i;����є̂AK� �Ba�������M�l_�˵&J�ޙK_�Oz�cH7����� �J7�vY��%�����j���)�Rb��F�$	<GG|���{�T?3A3%���~�#����;�;�Iw\��:�]��g��������C#�6>�b�rB�8��B(C��K���r��@OS�2'􏕌�a��y�7�����*8�;?�3��P�D���{喝��z�vc2 t��+��%��}8j�3˿?����Bm�'�fi�ñT�|��R�;P;=�1�Y�LLsw��)�aԔY7_�M�7"?i���a8��ݥr��ePL�O��]Ye�%K?3�*�o'�ڸ2m; �P�r.:x��~�-J�	�P~��XB�%KH!;����U�u% 
�m����(d�Jk�	>��_�������{�S���ş��ɚвV��d��;*�+mH�������6��EB>"P�K(����)�
�����Y����5����F��z���F	�V40�y��"�����x6���-e9AM�A{����!y�R6�h`�ȯ��	������s�پ���0)2���[���&H;��A�)ur�~*S��ߦ�G�x�muK�X���ߨ���и��z�g-��!���>��aqIn���6�V���#1�O<��<Uʆ��3o��tF��W'߃� .A}�Mw��|�kK� �	0�X�����I����kXn؋F�v�g�l����Yl�З��"� ���zC����	YY�Ik���YY�|���~Mw�3�'�&s����l��;����{_�F�--�鑹uiV���/\w�ia�0�M�Ϛǰ���_�dߊ�9���.ҹҔ?�=�[00���3�9�Z�#��MYM�$�-F�%A�d:�c& d
h�����^]�\��bG�@���C�*�Ïߏt�QII5-��J7ޑZgf�B+��L6A�2��ycE�T�+ڦ��cyl^��Xd���7=|����v��d!������ \��v��(t¶�����~�9��ӷU�ń��Q/����n/��'�B���$ �]U�bM#�N������$vq)����3��
1"BRXiK�Z�Г��_���M����h5���C�{:P/��c��M����U9���3�����d�c##�ċno%� �u���cf�������v��[gF�:Y��U��?��]��!id!�k��!G��[	|�^��I�wZ� 5
�9�6Y��%/��f^�rG���Lkt�@�':�#��=�y�C�%g��c�sv�E%1U�9�׼uС8�4�]�!���
(��B��M�rV�dw'��Qꂋ��gt�RQ� � �Sz���d�r'53%�,(|r$��!����ߍl�	�F�]�Xr(Z��""�IS���y�o��v�,�צt?�iĶ硹��hlb�EQ�ؒ4���͓���%j�m��� �n�#=U�CZ�mB=�%�W"�O�ZH[�{ЁK۬J��!���+"�FP��{�_����hգ�}�Q��d�1� G����yvHtpN�7�O���**؎-ח-� ��@.,`
P2e���"~5�LR�:]�_�׉%�?�ȫ��g��Þ���T]�.�����>@` �"�D�wѧ��i�"��36#��e{�&^����%�(}l���,�v/��C���.s�4���ѿ�r�Db[��z8}Ѱ���cBDY��+6@���j�;Z�itU��Y�������f�}��1���W�7��P��4;!�`A9����@��@���ڵ�;�.�;A�����	2�e�>��|W�p,���鹵tűJ���N��R��ظ��H�@�uz�A�ǒ��h#țџȳ�s��^�Q�x*�5���n~b��X�7;в���Փ�_�$�u�׷J��
螓o�Y�xG��r�k�B̧>�u[o#
�:�y��C+�����9�o�֟���obVTD̺�����Ys�@�����μ��Y�>}l]�5��b_�j���T����y2O���	���d��`.`��\��c��{"�Cס\�Lqo�(�����pW�k�����@��ҿ�l0��5�박~Ԅ�B��m����;)XF�0�OT��s��R��7������XI���ʲ�r}���"#��Rԥ�5ZgrI��s�]�R�z�Z��ȫ�9b~,	1��[Ôi!!�,�REw6+7�%YY���*8�1N0O�+6��I�iPE)�Rۺ��C.y��(�� ��.�C������%�B�zT�F&�mx,�S�Q%DI�p��%iE(���[?H��z�^���:-@�����\��$�~�εy��B�����#2r�I��%(2�-	ʢ!5�=��3�X�d�/��Rc��E=lR����(b�T��`�ڙZ�f�F%{��ILW�`�*�~�f��h���T�a����V��~TvOV��ӬCl �pn�M���_q(Cz�"gb��z�FY�S�����Ľ�a�j�
Fy{�ӳ1����+�ﾝ��1!K7�
�)�$����E(D��6�d߯�4le�|[��j%�9�͟����/C.� -u�m�]<ג*j+ɳ1I*��i1�+/6Hf5_����PL?��,���=�Z�0~�u�R���r��1�(¼c	?��'�#?� (�Jdi-4��SO��!}�U,7��,�^�;��1�����a�{�O�PA�/QS��́v2�ٰ����N-=Z$v�~�= 5�7|f���yA��;�K}t�àؿn�l6�y���n�aCϞ�XȱynJ��j���j�n��y�P�Ux�/Jc�9��pJط�|E�ަ�[�ꈙ,�!�?g�ˑ�T�j �[%�l��`<|+�,z��{b�*T|b�o�μ�_�CX��EO�udO���._h��@sc}���r�
���l��W}���uU�b���?<#�CNZ���h�Z��we�S�	A��I�Rl�F+��aF'Q�G�K³T*�^�ݚ�J/���bsn=LQI��=97�S��F�N�q��Ύ/�B[�p�ـ~��C�O� �cn�;��`�>�ɧw ��U�/���}����J���P�������۞ؘ����}���8���~!����zSB�@�n�8#�N�3o3��"PF.򭖵e��_�&.�V�P�v�<C��K$k3������ج��?2J���xz��
b��g\�~f[�j剮�+/sg�3)k�7�럟lba��,�WwC0o�n�QU��]��s�G��""c�	�N�:l)�(����jVe���٘���~d7�Y��8�:����t�S4�g����ċ��耶K*PT��(����O'���p�i�`��J?��bGdXr�K;
C�aӪ�C�<C�J�K��RruŊqܻ�wH��w]H��z �Q�����`G��Uy�렽�5x��E�}2<�Y�i9�DQF˲o],��9�!����c�i��j`>.�������`�A�񎕩l��Wa�-���
�Dq�	�r�`�,C= se<j�k����D�2����N]�V<'�5�����Ô��#�_F�؟��f-�g��+@�kL���=��oO����$���ybȆ8��G����g��9�0v$��N#�7�:��~���!>Y�da� �mwU	�5�N�k.f��h�R˝� A���JſCY��>�M䟎h* $B&��1��ZfOhv=qC��P>���0��{|�_��������f�����	��-�.�t錅��C�L0�8�/c��;ΎV�qך��M���Ȍs\#u1��ͮ�}c��ON����[,�O�yտ�v�#��D$zx���$�Qh~��x�����Ŵ�k:��G���B��ِ��|J�}.�$u|ɔ�J����;=\)�|o��OѤɧv��}cXM^|;��� �o�0T�mEC��D���s�Ϭͼ�a ^x����{�岏�.��,@�m]�N��E�z��I�����Rߘ�@c�T�!*6h�B_��SK�^�A�Y￳�T�9'����r�I����sÁ5��$YkA�z�������8��T%�3MV*���Ky�8Y�O������^�>75״c��<t8)���eg' ��>�ȳ��|�P!EB�P�����%�����"z,\Uq!��-�4���:u5uu�i1�.�Ъ�6,� ��?8�t��$�Z+L .��x"ƠlD��A�h��� �NgpK���1��#�����1P��fN�$}��4���7����_(��!<B�n:Ĺ���9P���������6��DИ6p\�<�F����ů��zUa��w���B2a�xP�!qJ�m�\�,��Ԍ����74���\(��9;�x�#��m�S�e�����Ssi8������hy�a͛�=˭����z���e�'�Ӱ=8�đs46/yg�qF�h!f�pG;��4�85�?<�fa���G���ߌ�9Q�k�����A�� N�x�F�x�YH�F[v� 鋬��v�=�����5��K:X�1�ϟ|�J��L�	h�ZF'm��8�+�����z�?�+� ��~}a���3�����v����O�-�%!�1B�@ཾ���l�K���qG&~s�l�om�����d�'g���6��愦)DsI�I
�N��N�(Y����V��IN�E��y��E#�pn��>�7
1\u�]bz�n7�/��]�[�Ѿ�O�m��)�|x�S:{�W�s��
���Lr��:��H�����тaLɡ:�C���IA��;���0Gd}A9�(��7��5r�\��D����iMtL]�PW�qыD�9;�_p��b;��XP��9c��7hM`��m�l瞺�٩������}�+g������4�6L�3r FMǚ
��Y]�4�ݡ���<��f|<!�W��?!5�I����� m��ٰ���T(�ǛJ���i)�Em��U������U|y����Q��Ԛ֚�h�u�T�1�!l=�JE�3L8�ɻ�I��a��,�5��ѣ���k���0��
.���,��P:v�I*�I��Y��E�y�7�Hvd�	a�
�������Kr4�}w�bǨ0<?�q���*���`��w�r���@5I�v�q���&�m�+�m-�o�vO?�L��@f����e�0-��Q����2t�M}�����5l��2oa�����e�}~�	���(t��\�/�bz�1ۋY��܈=]�B}��D�j�X�Qԥ��9�MD�S�A�K�B���hFۉ�v����r�#�b�R�.�RT#=�jk t"�WFiϬ��א�O���W�+Tm��f�k��O8��.�[���T�`�Z����bg���_�����閧ZP���X&�|C���cl{��ɺࡶoZ,Cϵ�Ʈs|���/���TC&�n����nQr�s�Fǻ�m��<�O4@�>c�O�Uhy:����Q�ȵU���Y��
FW��,��
����.�������`��|/���评����B>�&��n����Ѓ7G�>q��mO�n�4��{���(!�ߐ�Pr�'���T��w��1oZ�	}��VJAZS�(8��L�^����]�A�4M�%8U(@f�SQm[���;�W��g��WD�e���dk�K�U���
'F����X�Ѐ8�No�?�9�pMz��)`����hT| �B��a:�:�>��|4~r�D��>�2g�W'q�E�I(~��t^�"��,r���@pq��w6|���FWȡ%*��zj-��im� �:4�J{��IlǷu�=���[N�_(Ѳ��>	��L� �DZ�2T�8���b��Ue]t�����]\�ob�GK�%.Ų���/\�^��U��ER�t�Zn����2�cǽb� 3�R�K��/�E���kR��)�_���Q�X�v�kXT��fl�wj���E/.�W;��E�AVe��~�>-��I�Y�c�cʏ��3��� �VU*XK�w��MK�LC��<XطxH�gL�͑���7* �eb%"�S���y�"+i��r`�E�d��6�8F_�Qݫ�ޟ�ʩ����"ʷ��z�R���T͊����EXZ�6�)�p�bN��L�	Y������|�QSw�����6��&���B9,�W�umX���/ұ�@R�Ֆ��X�
�E��X���H���})
��dA�e���=�x�?����ܙ�]��`�\_h0ᕱ��]�W�X�~�H9r�5�� ���`�t{h��M���~5���c��/6�G�eƫ��n��`�~��qĮ�-Y����fO��_�1�y�%��7.̄��;��҆������o�5��#��f%6gG��u#�u)W�'��$�[.��y.StVx���4��1D�p�og�����
��%�]�Ll�YM�?F�Jh`L\rP��1���Ӊ�Wj
�,;U�Z��O�ԫC{��Pŉy�m7i�6	�H��a�vPH�4U8�v��B�b�.�F>&�e6�A���V�[9rP<4׾���Xkl�y�Wѹ�s�9��d`yL�1��肂S��낗�+�>1� �lj���h�6KPn���Bq:�.�(J�3%7f��s��a�`j؍�E�_�(�}��2A�7s�n�ԒG��f����n�Q�)��L��%�G_�S�����b���g��GU& ��˿�5�T��@[{M�H��H�C2vp�����Sׯ��]`	5�dk/�0	*�;��4��ro���>`|w�ww��S���_&��IM-���]��[R��e�Wr�ْ��+�`��}�tu�ڏ�d��H�d�l�ե�: ����l;��t$�9Q	���]����C=�/e���|�-�9�p�da���[!=��ZB��4�U�����0t���0ymG��ٓ�d[ۑ�E������v)Ҁ�� �G�5ndimn]���b��1�
���x�տP�x�^��ts|��f�O�P��n|�|Zl�n�tuR��YG&2gʌ	2��3�!�1Y�z1����O{'Zq���5��O���J�y�Y�2���!1\|(!BՕ_�s.e�AV@2%�A�;���v��|�r��.��|$����ʬ� 3+�z)p�̼uh�ۅ"��l���$}y�&8�B��!aG�F�6 ������è�e�"0"��_q�Ɏ�?H���:T��(��y�o�{Up��I����IG�2��,byI�/-8�q�.���U�ڙ���b]ض�����6��}
�?��?�v�@W���$�_�(�P��6fC���3o��Ŗ�a�ֻ��u�f�߂�K�5㑂�ܑ�nD�3PT5�F�����!
d��*�������74!��~��] ���r���� e�j{���7��ا.!<���\�6KѺdp/_/�q��yD7�Zwo��^+FJ�����?5���$w8I(7�Y�Ȏ	���>c�d�yJ�d���ج��0##N�C�Wb��K�B�o�q8��j@@�#��6��pYOL9m�J�E}�Ǜ;@�GC9��GSaLک��.��!$=J�}��k�O����~l
m���5����vj���Db�{J��"����T6�c����6�ò���w�a9��"��_�ٯ����L�v��+_4�6�fV��M)w�+�����Q#��_J^)�S9���T%��q�`D��`�/@0�kv\XZ�#��#�����_��!H�c(����3J�{�S�b���[y���ր����u��TV��K�`b@���p�,�]]��悷LqC>%U��[T�W��=����(��c��>-�9�C����o.Fmq����@�H���z����-YM�ޮ�xmhǜ$�m���*�X�,dY��VaJm8EuH8�ˌț}���l8,YI�v�q&!�*�o�_8�^���)��2��k���������̢�A:I\����9�c:�f��O�['Ͻ��������6[�9�:8����i7�j��u�b�����IM��~��\�Ec�~�&?�켽Reb����9!�&�G��f�Fk}�o�Mr6�eґ��h�u]])S�
�\8Px�T=ލ��z�r5�&k�/����DKji@�ᤃ$�x�J��M�-��Q�q�l�����iJ��C2,stP�`�I��?`h)���}N; ^��"�l�������kC	�(�������D���p�+���q�T��H��ܾ�ox�lq�'�me�M�*h@������|p�h4@:_�93��@G-g��;��1`χBg9Ƣ��9��o��(���&��D��X�p��b{m�p��z��(:�U+�qJ�{D�S����Gf�a�m�D�9�n�#�~�2�z��0P����/c%�Ƹ��6٤8;��\5�1 ~I+�K��Z\�n�`�vvy�C{m�=H��)�m�yBy�N�����h>���Ib���YS���1��Ew*Ҝ��N��U��O"4���M����a��i'���E]���~�`�8��>b#��K� p���l>nJ�	Q�������X�8s,���w��3�U[�/����U���+*B2����]2����g'u'.:�ȚlRe�ο��3���Lq
b}?r�2���+{v���,��?%�8�ʇ��r��[��9Dt��Gr;������9|�\�t]��hn̪�_ZC�y�%��pf�=�
P��m�s��7�&؄�!�ʤ��ϱ� <�Z�Σ�pް��/`�(͖pv���:�����ѶϹ�6�V�Μ�ӂ��zꝘvS�Ԫ�	uF�������ʊ�)��z���Rg~�v���F	�W��B^Y��r�n�px�寂������b{��ݕ�-��~�v<-b%�=fMW���$��^�g���*��=�R��<����*+<��e���pQ%��;���8��f���fa�n�V���޸�)��+�����[��:�Gv%4�ȁ�Oɭܲ�e���l����L�:(�y����tww��ط��v��ڰLkq|�	+�8H���v�_傢@ȩp�9��}���P�fbw�wNCL
L���%jl'�u��佂e���Z��ܙ�
x�)�c)���@ ���4�D�� ݳ�c�o�d��5r�t�8W�<��>���n��򐷧�M���E�2�Ƕ��O?5P%i�9g�+D*�H����-�4�_�z� ȇ� Y�e��!�:G��Su���\�R�N S���:p`!Ob��>L��Zy���ʩ��k�Sj���姴��y$Ufz�Dir�[NNV�8ߟA�W���A�o'}W�|U�"q*������>�&]N�F���ɲ��ה��4�؇�x��!#4TI��`Ō;����up!h�hT"GJl;�v8��-� ����~�a�Zs����|��.N`�V��K�4ɸ������u� ����ل++�+(=)�L�o;��g9~f�*��i�+(���S�$�f�T��6	@e���C��*�Mj��i~G��?��ÐN4�Y�e��O�5�?�ƃqAe� y}}��}�'��6�f��=�BްO��ݿo���+�ؘ
���F�7�=�O��4�Mrp���I�@؁�B���aX�xᾖ���hv� T&j�zxY_�|��� �`M�Gډ!�+b(ec��)6���� 7����!4�2�E�y����Svq0�]{i���-3�ҽp�$�
U{-���ޙl�N2��J����j��8�;���t�Fq�rB"9ήoV��TdV����Ыy�[�<|��TgO8���!���9di��s`2oc�4:�7�H�q��8Fb	� OQ'�Q �����^�x�Y�������3��+:�;�4���#Ï�7�\h�XwĎ��|�%���0MM����3�aH/�lW�g����oM���0`==Z:O�����L5��P��0]h�i��؂�׬�_O��Gkn�������z����{"�o�h))�l5)+3l��3Ac���D��=Omݜ��́�!e�L���Ę�U ?󅟭�ܯ���ũM�~��	!Mi.�S��F����AR�V����i[��m�z�;�u���펚� �J>a�v�c��S�O��Ɣ�IZlY�����^m�?��m�
�(�Pܖ��z6�Z�g�!��������A׾tWB����d�ݑ{�>RN�=��&�?��WH�l�����od��[;5Ha��6�U9�2ګ�E6��C�h���o��5�ϲU�i�[/.j&����P�V�������e��Z�U�9�5P��E��G���k=�c���eu��N풌�'�v����������Lʈ�$^�n����'F�6@�tyH(4����"y�<��;UE~�q�ۗ"�X9�3�� j�C6��T����29bj��D���|7ͨZ �%�˨���R	7<Z��bX|2zJꁅ]\^G]�>��I�C���T���b{x=�Je�ֽ�t��l,�v�=��l�>� \��A�OǓq�n�o�6H�Ⱦ��S߼�
"���t���9���!3�ǩ�/+lZM&�
�33(ϰ�Ҁ���,����Wz>y:��=�~���n� R֮;�y���K��Y�]q�C?c����Fu׶V�#W�ܧ�
��π��H�E3c�	?3a
ν��1�{����'�}6��;(���Z�=�y*!�_vU�%6��b���"�jBS+���D6�pu��V�����Rn�)wvJSG)r�a��̛^d�H�X�t4HH\�ܺ��x�d{X8u׻��a��lM�8���XlxV64EB    fa00    2730�O�$.��<2R�������zg?2�V`��}���mn\�>#�?���%�N���,)���6i��p���p,�yj��s/VI+DT�[�~��I6Z�k�LQ���H���<%�~�����Y�	|&Z��}	h����F�4		l�Sh�x�L��\�����	�<���V����=I�Td���Y9�=�P���d�����z�Q�ubVL+��b}"X�Z;��M����	�.9�?1==�~`8�����8�g>��;6v�Cw��Zd?�w������Iu4s;I`�\m��1.@)�7]�D'����J���x�q;	`�C$W>8zLi4�� [���t�b����.~r����l���p���pǅ-��+@:}I�1cP�+�����R۫"IAB�|.�I�r��_N�?p��'t�A�}5�'�)�ޔPR��S�'N�����_aa|�j���!�{�&�f��2	��O�&u�0�ź��xR� V�-��P`�u���* ���A�p\�-B��]6,;��J>�4�-��\_	+��$�oܻ��}qT T�`�f*�>^W9��kq�d^�s��pV�˱�"��}}%�9�+�{���WV�UC�=��Ө.$���tQ\�;T�G�f�Ҳ�u!���4R!	��7Gȵ�%v��+Oj�w\���h�0'Gpdj�nn�t�Б*L4Qd�z4ub�hϹk�4��;
ݧ3�[���"Kj���n����^*=���D�(F��=��?~�g�)FS/�o0�@p�c��ϛP������3��n��^�P�A�>-����gg軒c}Dȉ�]�@�,a�PUv(o�w���r!q&��'��TX��Y����9w|���&?2�$�KuT���t�q�d�@�#vjy��qٕX���������ѷ�0i!	��ۣl��4+���LQY�(sXފ�3��y��X~�A����h=m��Xک���(]�7��p��Y�˾�S!�D�9oCN����b�Ww.�d�j��2������*�W�A'��ڞC�+,�G_��q�!��ț�Cɸm��n~���K��m�W�B-�m��C[ք����&!�������Hj0I��p�T�]�q�v���bì���M�x�le㽓���$I^���$�ݮ�O��~��7>�ĩ�k��o�IS�p��n�Q��練=���'e��.ρ�'U���Z�O���K����y!�c�W������7uC���
�ȻgȍGNe�q�a_l�lQ3��%j�`e��T��KL�߆Z&�	}�ŀ�� ��x�������<�|p}�Fe�Ck��. k�%���l�'���*P _{�5&�������L	>��\O�H}�tv1Np���3̑��z�퍢g�"nV��[�Sp���*ͺo�&ROIW�Ά��qJ��:4��wN�A��N���aϞl(�:��|ya�i jC��VН�0zё@�9��G%��sLZ�c»�O�&���1�/o��Ρ�v����b%BL��B��P�_%.6��Z�������9����"H����#�*�nN<��x�A���� ��KA%	��(�V������Yy��R�6^1�S���s��t��?��Ag������'���F��^�A��X,�yu?Ҩ��C�Ճxm/05���8;�QTXQ"M	$���[�E�͑>'ӌ�jāZ������QO�\�h�~V� �4�@�tn���Q�=�%i� �U�'��%3�8�H����'���Q'�::2H؍K�-���wTV�{���q�8�5�W�j��n�L�;�^j:k�[��'��<�֡�,�?�q*� D�*޸��EFJ���	�� ̙�{/��+�6(�d�Yt�'yy���C2BL2̈́"���z�����&���^i��+�~�����qm�*���m�'�����]Ϧa�t�[��t � fX ߣ#�_5,��4msϠ��%`�t?ȻmЇ�U�LٵJ.uoZ@Qy�㓟t~��� o+���&��nZ��Y�� 	����σ�[qp�������燜�o	��a}���%ڧ#j=���8��-$����
?�5F�y]Ͽ�F��@��n�~�8���}�� ?M�b��YCq/�����{(q��Ew�38��=���#[Y\�8��|���p�6Ճ-�wRl�ppkS�?�w���K�t#qۮ�f��.�4�+9:�@V�<�%ABHzQ�d"�k�m-g <`�e�(6�vLl	�+�Z�A��C2�y���@鼎.Z������.i6J��&D�W��l��a2�
$�|Nh	̔�����ţ��}ZJ�VMZU��/�K��ќ#�֝�nK�ˁ7%+���1x������%��3��j�ʢ�5��v�0���*��I���k)@\21�!�����i�������튺f��'(�E*��%���dTb��T���Cɥ9F����h�ԑ� 4�S�|
=R���T����!� �6K~��~��3ҠW%*f��휨q+4ӳ�~nm��ma�YiF��\��jq��cHt��ͣ��
i��E8Z�ΊW�g�����<(�&Z8��V�M!�b�ѕ�(�.s@�������ʵC�ӇvO������7X ���ӭ!k�gί;���^b�'#�%��88�����&iԭ=�c��6�����9�@� KnQ���F���
&VV0�#��9�z�w���
�a���n�j��y�͡��̤�n!~�V�	Q:�bċ��Qd���
��!�hY��O��\!,d/9a��'Μ�w���<�ԍ�����P����:��k� �/rVdQ�cKj���?Ӏ~������2��u��p���Wvѣּ/ǳ�6'r��]h+8^i�S<����h�^i�/���m�1+D���\n���<����4VᘟB�5�� ���ǥo�=C�~,�y
&�XUw&�`V�X���].��Wq��Q���.�t�Q�Bn�u�9��A4π���/f/��~{����)@i��-��6���֫�a-��_�}��~Z�:�w6S+���]P�����l���;Z�oU��F�O�Γ#�;c9	�#�w�֬=�ӭ��IQSs�����-���U��%"Qs����2	|I�ٹ��!�m�g^����v�f�,�rؐ���� ����8bҞ��(���U�}�6�&�ޚ�aƲ�9#Z���L�x�Զ8��#�i�S�T��:�2u�����2�u�	h��j틅O��I��.`�I��[�f�#��>]�	��<7��e�A�c�u-�î'�k�!�������m�'V��Hb����'!ji�!S�%t���)>6g-�+s}�1Γ�~���G��q��MgP��C>}Tls����0�$@���\�@�ؠ�g�,n�/��i��}�^{���s]��5-�ȡ�&�b^~�栲EL]+:�)Q�]��O�Y�d{�z�����w�+S���P����Չ��dJ����OZ7��+ke����H�_Ayn*(��_���%n��En��|G`I��+L�/}��;
q�`�J�W�w8��6���JC�(���Q���f��ź2f��."�5ij^&�����L7?�C©a�r�a�c�(�Q& �28���Z��o�X�{ܧ�W����uL���֚2|�v@� ���؟ֆ��e��қ��JJ�R�#�nIt��>4͓��Ż'��gH	�B���Z��x�\��U`�ٛ����竃���QZko��+��r��F'�mf]ꌚ�W�~��8�V)�j�7f�6hYWX(^�|�zC����4n�c�}U�%{��4��q3�<򶊻���0��Zs����cN�h>fۺ���|�0������q�,����q����l2Z3���(#��W���y�`�2evu�O%ӆ�n��LR�gm��T�)~���G\��٣sI��j�\�q�t̗�R�]���ډ����Q��{m��O�U�S��縰�F�K� 0��e�)�������p6��8�J�[M�]#�B�?)�|����%��:���;֪����_�F�隋MLͦ�_0���P�q�Sz F��4�Y}�e�R�%,�A�p�� �:��6O�^B�w>[�ߚ%A��I��3�_(0�Q7(J��l�P�����ߟx��E�1C*]-Y?��>�q@E0=+3�ѯ��w��k���X����0'��
Ω��ȭ䢱&��U��'Ӌu�sO弐x4�DX�����K����,���A�?�c�x'���x�&�6	����QR�u[� 7��~�� #Z����UA�R��)�(��G���<��'����s�<�Y��</��S[�'��:L���[t�{ê�Gg�D��?H�Y��R�'@�+��;���m��x�F����6�3H��!aj��Q|�ξZ_l�(oE	)8|��\�5��].�cx�����&y��薚WբHe��U��2w�jht
�ί/ϳ�>�!O��`᝶��褛k�Q�n���U�����M�6{4X� ��G����&"\������"������2��'�7���� ��_/M�8���L�"ozp��eO�?m�!�bL���l�'o�V(��t�^�n�C#{�Db�h�j&n8͐_����ֻ,�ed�����C W��x�:|pr������`Q3a�@(u��,uE#Q�O��A5��j
���F�P2Z).���p�J���ċ"�s�I`2���p�E8�CG�/���շZ^����g(�[�t�zm����0�T����~"���ۑg��.b��%8����M>_B����"؃�T��������Z5�������z�0`l	��&D~��Ԑ�웬w
=JA3/�6���Aʒ��ϓ�l����g�*��gwu�A�V�^������Q�7EX�y�	��\����75/֏�*o�w�ȵ��a7WS�TJQYy�.,c�B�<i�f�2ct��T0ǀ��|oe1v�ӅM@��"��좿ڨ�BV=�ᤗ+�`gg����F}m�p{���S�e�Q�VIe�jV��t�)���)@Y��Fϸ�6���G�<6�C�1���(� �)��%|����<ϯ ����҇q���B�����;��7Cf���mv�oTm��M�	������.���0'o��z�1�R2H�1�˼�������5N�%��y{F�QE���:Wc =p�:V�Y�T��9qx�'jK�Ƚ��g�,���m�����x̀s �W��L���h �J�e*	�v�,\���'*�,�jie��~ѳ�E ���ػSv�:��+���#=X��3�7�q��0�܎Vћ��Y�F�?�!AD�S�"1.�Pr`��;�/����Tf-=�ɟ-���{��h[ǄVpZ|���Ēo@#�w�(��_�*�٩Kbw������Mw��(}tU�&�l��W�.��tt�\�UW1��Mr/p��ច7����?��A��YqV�GY��GC���%FR��N{&G�qy����8�# V��u\H}�,ŮX.���;�W�:m��)r��T0�+�:�T�=	�����Ԝ�O
#~��rR�Nk������Q�ì����Ȥ�;�!��Nh�٥q<_���8I�L���Q���<�(o?/v����1�D�*���K"M�M�KZM��-��9</�m�,`1��B�E[YbZ�a���0������[�쬷�E����o���t����ښ,O�ЌԀ/����~�im����Z%��.�D���X��X������u�S��@�&��8�u��x���ܪYT�T��W�Z<;�[ghF$13��˵|	
m����Rp}�J����
Zܒ�a�� �Ж/"�dA6�`�^��s�C1Dv�r�I"�w�O��y�)��J��ii.I�K�*���W��G�Ɇ�֎z<�)�A�"^���:�(��=��]̿��}���8;�{��c��@A��g�B����uVt�V%���W��e�^�����7�)�?ߣGk�{@t[_Z�WVe
�ϥ���,�LI��A���;�ϵ�IB��:�7��{�rܲ�!O0���9���b� �����}	�.1�
ل��U�.	����t��d��6���=\4]LF�ݝ�}��������3r��.z�m\o+�Η[@���ZZ�����T#�{E��N���Q,2��� ��K|��(��Hw.I��/HJ��1}��V]q��Ţ�
sB��4�!D�25�?��g�1�W���gLIH�[��������%�p���
{�c�s����5b붆��4IV��#�������ȗ"90����B�	�Ve�+�`s�������5	5�-L���O��w���`�:�8�6�"�B��u�̜���h�uEg߮��N�͖΁/p1�?;��]Y__:��U�in������������^UO]�fA�L\�I��ƙ�c,��H��{�2�H'�(�u� �`�[�٩Z��JTPAn�M95kk?[kf+u���=�������������v3�+W�O��X���-�!�Qr`�����Y��\ Q��c�x�����b2����=ǬW`2��P	f�]�`�@�4���̏��E@�$�}�Mq�`s�4�%�G%���	Y4?گ�dǃk\���O�J�ԥYA M΄G����^^�@����Ə���0VE���Bo~q��e�7|�F�B��2	U�量��1E+{G��/�2����i�sď	�II�7�u�)� S�> Um�D{�ъ�rV��'�,D�@�]�4 X�c�[A�`\��x� IU@A�U2n�;(0�s�#�[J��wl��ߘd��Ñ��y@Ȯ�K^�x��-�=�ZsXz��č��>�fSgg[ď��Dʴ��Z����\����0��jq�̬>B�qiy{�g�RS��Q�ӔIRa?KZ Ƭ�ky��~��`����	\�GI������Ak�
'�C�u��t�#\��
�ǝS����P�;����F�6H�)s�)w֩�<�S��ʭ�ȝiR�
�h�ʄ�rhm�x�^��W<P�ʥ϶��PϥaYg[	al��1���k)��\�	�
5P�KV��E�u.|��'^,}�����Y��I:0�� v�>z&�q!�j�!p��&�[�^Q�A�α��&ҭ��X~3)�'��ê U�PD��@�V�0�\�t�}��Ƣ���D؂�ķK�\~�w=�M�	i���f����G6A����GʤF����l��/�����O{T�XQx#�P�w�l�TR��x�Q���
pw�12�?����6E�϶����0�������,�=N��W��#��ʻ\!��Z���@�h5Ϟ���:�5a��pz�w,CIn��<�,.�=��B\��A_���1Ձsy��{�����Q�1�N�1)Aqx�*G�¤��RD�ӆB�cqS*����6*�*<ޮ�z��3�}q*�Ś7[�X�o�HD�|��M��q-z&ޚ�3
�Q��-������rf�Ε8�����s[Y.�#���*3�ťn�^ۺb��TSp�+(�x7�\���+4��Z��Z9�H��-��(b�^��S-V�m`� ���?�sN�Wv��]�g���S��Ě���̯ P��3�W���~}�VW��mJ�!]u�����c�&�:�T1p��s�I�������A(�s�+.��븟�1� �H��i�DP�VU:V�L��C�U�qˊZ�D��SN�X��&$�j�uPRHu=7-��� �.��le��^��=c��6�(IX�7V�-cE�H�4?���z� ���(��~\���N�����΄N����j�����~A���F��ɕ8�Z֊�y�Y�PEP�(�B[�{g��y�����--`�	��"b�����8�P����^�Ą3�W�E�<c����S�s��zS��φ��6�=Qs��֞�7ĩ2XT�Jy�v�Ad?�`<���΍�c����56��}���8�@E���>ލDH��l)	q#I�M5C�$���g��=�- >g�����L:~A��B�Fƌrc���,��1br�M����V��oU����� ����#T|6?�?���mJr���� ��N���q}$uX���k�#.�y�$p���{�I׍�����kBS���lw��:��GY\9v�J�w�Cj�W;����9�ڭt� �%��>H���N�9����Œ�5�NTb~��'?����B6�;%�_�L�L�F-��d�)��- 6Jf�,�mN��DaKl������-�Y� � �����
8�s�S��֪�Y����@��9��xӖ���_�@r_ak���p�ҙ ��h������{ק$��4���5y~J��b�c�;0 -���3:�/fe��k/h` S�i�*>� ֩�E�vt� I�,�G�j�-�P5z/���}!HK,lR��	4�mB��L��&�39�����Y��3�C?m�;w+{$^�}��%���.���q�c%����0h5�L=E������S�l��E�����~I��@�l�����u���R� ��0�g��p-�2�%6�_���f����c�pt��݉V<�
{�B��"����'H��l(��H}#2CR��P�d��B�l�"�C����F����Aq~�!`�z�l[ 6���k�S�Аl��T�@�B�U�M�[���=M�i��\O��)����N�0�F�a�g-D�<�8%Y��fs4�!@$_���r')��`��@���rjёE;��F��{�TT�G��.�)���t��>5���aB��-#z���[T��s��w��ta�Z�<B�!�f�L	��ij&�\�9��)�J����K�
��S�Eܜ��:��#^�V���*���z�:׀@g���~񉚻�;�ˮ*�(1lE$ 晙闱����1��E�e=>��]]�	���!�Ԧ	��RUT���J�j�8U8�~�v��`x��D�hX����n+2�5�zV��YuRn�����[��;��}���ںtHֹ2h	")��\��2�!����`���flN/6�`#���{Y�>���QuJm��+HMD�N���&A[?=����t�K2��	�_��I-���1z7��v�c,n��t��{���4YjeI{���e5i�
Ȧ �
�lc{�R�O��ac� ɥ&�1״���&�E2��W�Xbx^wQ�c��f�L�G�Z��X��g?D�" ����v�O]11ā9l��I�Hv�(Z�GW A�m�E�^oCr�Sc@�zY?����w�����rhY �-	�
���U'�x�r���y�@�T}("f-���4F�#�8W��ϚuR>����-���
��G��ot'~Z0"���NK��G���畱ѓ����w�W��U�E�M�jL�����,�` ]iD2��"�I�2.^7�9��ef�_'*D�?�՗tז=O���6e�Ƶ��÷���x����sv��?F�I��2rj��T�s���gJg{R���������P�/a¿9t��'j��K�,�yz�
�lp2�J��$�ʫ��0GL��ۭ��O��	�2C�[
������4�aD�����ϝ��O� ����ema���=�$K��������+s���cM�;^�t,Mc��Dc���2��60,y�'������`x��Hӂ�\n:{҂�3����:��b2�WV�ᦑ�K.3��@��a�<WUIy�Rv�Y�P�GR���IU(G!�����H����ζ]���mנ ۢ��6hl���}/H&�����c���P�����Sz�l�Z�� M-Q�A�8�XlxV64EB    6356    1000��B��ͬ���鬋j��C�L����6�4��f�� v�_
`C��b�!|ϡ�Kxm�[*�����&�M	�'Bk�"~�l�)����w�+{۷�V��U*������@ߩ�(s��}�� e@��Չi��k"��>� �R)��l�@�V/sd*:�T�*x������r�1Zh����q�[��Ib��V��&ӝ�h�ҁ�&�y�M�~gg1�N����'M�-c�U�E���/n�g�S�_4�\��!��L I��E��h�VP�4�W��2�tU�2$>�[J��Ή}�g:.7ߝ[:	�����qIv�H���:�8�,C�G���f��"6W#��B�����I�?�H��+��+�;��+�R�,}�R@*��4��c9�d(td�	�u�׿s-��ɧ_����Zk��e�P:�ī����VN�iY�M�_���9��-LGP8�b���8�˱�Leor�-��=�&�� ��2�ڪ ��l+�!j6)@����V趾�|��� JCHH�叐/��-�����7(}w��V�Cg�J�:3E18���EW��D��5���S������VϠf���2�M�ȮP�f��Z.מ��;��IL���K�n���ݲ'i�|�����0m� �� �h�Z���Hڨ��6��
XE���kc��l�J"dZ����J2���\�c�yV<�|2Y�IԂ�'�t����W�U@�=JS����A��aXm�S|�D����n�s��,�)�0�/�z�x���h��;ڑ]0��7��ð̿������.;Z���x�N�-��6qyWd;��hp�+J���ݭ�?�cn����K�=�-�,�}��(��S��EC�.�n�~�N�>⩘���ˍCo]�l�YKiX7Tl.���Z��FOz3@���sR� PF���."�U����qG5/��ā��7����'00'jLٗj��d�t���o�(�e�gՍ�,O��lr�����K���g��Z��̃3�t�/�ҵw�e���N���\lX���O.�=E�i�9�勓��"�?�GQx$�NN� !�����M�J^Z
p��A��vۛ�ҳk;o��I򃆇�:��t�����C�t��@DPn�z�r[׶�sc-O�C�z!c�2y���A9��W�8v�Bh\�_Wv���# ִԒ&a�m�#pFX���QS]hn�(Ǯ�!3c���WϞ�l���!Bz�踔.�Ոc�]�R�Է�4ҥ��,0f�Gʲe�j u��p�E/���e�ct��@��fU��1fun���n~n���5W�������N�9��M��G=Y9B�w�IS\�I=�vΒ�;`G��]��9��s�{��O.�e�"�_�����!������� ��7�8r�	�A.y��ہ��$���Q[|h$6�l:�ī�D��=(tB{�Y��>e>gH�!��A���>��2,:t�.�Z�tg�di�9�>t�/"Q�F�QFP��g��u������ctx�� ���S6/jg�������:��&����$�&���n�UiD������/�߭-���y�v��^X�����X��`%#�Du�V�I	��o��=�l�8x��x�?��5�<�����Y��ҁ|n
T NjQ�|��F!�ðe�� ��T4��\�6�bu�WguSzjϼ��;{�'OCZ.~CLZ��c����������5U�}�Jg;��[��^W�&R��fn0Q?���p��G��@���l1/U8���:���C>(\ҊŁ��Y���_)�z�A��i%�hݑ=29��Æ�A8�1R��Ki|ߊ`�3�@���`���E�=9�ݏ�e뽶�:;_�y
-�.�y��L(?9����r	+~dR� �E�7�1����I�*�￬��偍
Mn�kW��W?���L	N%:�|J7P}K�7�a2�~�c-��r!jz�f⺆�k�J��bB?�8N�H��<��|�i�p���3��q�ofZWP��[�5a�����6D�a����z���MVit�G7~soR��	k�'i7���']������Y�����..;� ���^-�;�@>��]�w�z�9:�W�n���eW�Ŋ�;�o5�0v�L�%@�'d��b�:u^K��R2���5�o8�0���W�
穉��)��P��-�P��$�W��TMe��6}!.�|�퇿֬v/Z�͢
^U�*��#A�|!3�K�[G����tp7JMt�S�����{uD��Aw�D�)��I�V�zP��� ��Ū����u�bq���ziQ�ҚC�������r��
��dt�����u�)��{'��t�B��P���s�ϊ��*b�h��/9�"�p�KoPy��.����-�k�Hi������i^i�R�2;/�}�� �&��8'Vm�4p��M���&˔��̊Կ�Y��b.n�%�,'gy颍9ol���G�)�+./�I�h�;�P�bQ�~�q�yA�6*����Q�rX'�k�ܘ���E�H��ӏ�����F��|�08�ې(�K4 ��,�s�Ռ$�ͣ�j9)j�NT�m�k�4��-��7��閰>�z@E��r*K��Y]E��#�<�`P�&F ?Wlpx|�X��q��+*�Ș�ZfQ׽��'����?<)�A4�=%3;�����§7:����~k���9�p���ڂ��tN�{��׫*�%Mw�z��G����+O��uu�[d:$Y��r���e����g�����`�ܗ�w��b���
����NP[����=}�vȓ��uV�������:"Qh����r ��ן8!aF?8�bZB.��C:{NNL���W���s�~���X��[LŊ��hD.b��j��>O�*���'�Eq�7<P�^s@Uc��#���R����m}+�bB����d9����t
���K��+K��� �iNs7�s����)B~M0E�~a,"{��v#�)�l��_|�S���l��Ni@�| �d`�?jצYK����	E�}ӵ���▋
R���Žy�O��7����Gt�F��+Xk�B*7��1��p���^uT���*b���r�x�v��;�9�8��[K!��+B.��T�����-�x�VKQ.zz�G���'��|$���g)턲!�#�Z��`�.���!pU�,U�bKX�8�Csj�dB�0�.�EZ9T�*�5D����l_7_+}�� '
Ɨ�w�޷����H�N#�-�z֊ruRt����k�O\��Pػ	�:@e����'�-�����x�=��R��+C�ζ���j��v�Woʞ[�
�O�5	Ky�'�k��u�5 �ϐ���}�J�t��ş�����*��l�fL�@�gg�K�D�VB�~h ��;K���51Y�Z��4��H{�_)���<-���8�*ֺ��ZF���/�ΦIf_C�3�I��Ϳ�c����~����_��)��Y�4.P70@����r�_��+ ]�:ܶ��[@r+К�w��x�D����je<2��W�gx��Ȇ�$r�U~W7S����D�D����1v���ڣ��u����cj=9�xZO7�[UG`T����PMJ�4Y�@P�+H+�*��h:�U��Ѐ�Oo�3�$���1K!�?���ގx0�C���4�_�	B��U��Ux��l���k���a}ל����+^Q�A�U=�A}�Z��,��
�!�$������E�v�)�cC�~!�����]��y!v!ք��SX���l/&]:��+-	wV�OI���a5�PSV]|����m��^@�h:�@E0��^�Ű@�񦿇���w�ei�UBҩ���.����C���P�U�,�-<u�?|h���4^NҢ��
��|���aW����8�(Zw�4F�]�b�G};��r�v�-u�.�xb�.�m��l3��fӢ�d��k�R�膮+����F��4���ɪd`���HW��B�,�XP��Ji��f}S�=QʓqH~J����.o~C�up��0W�5�5X	������`