XlxV64EB    2a3e     c20E��YN�g�V�8m�����j�&r��jl~/'�2.]ߞ�TA��d��<� ���5�v?��������{P�m_���5�����4�0-�8����G����G����������ExF{�)�~/`J��m��B���g�����x����#3��G��w�"������)Z e��|�o�M.3�LЁ��	;�?x��l>$��!r
L)�bB�����1�|Lsu�#�-����XT�E�.ƽ:<M�sZA,q��f�\�<WD�(�:�YR^ax���tB%��m��@�Tdm��U:!<�k�o�<�܊OŪ�W��7v��̧��p��7�m���P����#�[����JŠE��Lb0;Ӻ<f6SXx���X-|՞�#6�vx�L�����K� !mZ��~��ukᔄE�p�������1$��4����9mZ�]��D5/4�.E����T��4�F�:��B�� >�b�ֈ'x ��Y�7N�������9�}E纺��c�Ɏm�!P�����Z6ޜ��K�����o��%��*�7B۾�E�h�M�w^(_��)��s���6�Qoa��׎�6>�ʹ�6Kb��?o
%R��ŵ�b*B2\7�N�Vf
f~��s��L�oA�e�
z���%��*��)��v[��L&�Z��K�YR�l��eg����g�F@b:Y's3	�S��	{�=�d�Xf��3�v��0�c��!��{Z�J ��pE�0�n��t��3I,X�Ҽה�S�a�(�
�Ol�.�nZ�Å
m��1йd��P]�
�͌pnf۠�%|`	�hky��[���m�&3��f�GN0�r����2��&���7�����EH�rv:����X�5础���O��s'�
�F$����O���H�G����#cZ�GZ��M�C��rQ���y��آ?��:w[ت�+mqo������h�t�.H������],zD:�镬�A�p+6|L*�|+vp����`�N����|b'@wh��qs���� ��6WG�0B
�pu��Dks��1�c�h�۽8ð���T�Z1�*�r�����K+��
�ز�F�MEo�s�u1i�&�5���-�JiGׅ`ud��k�;D=�Q^�ɲ}�@x��5�}��z��pQNz���w��v�+��K����
�
U�����b�B����<gr�PGI_�)� ̂�|ܦ8���V[��H�9���z1�S�֙g^�t�ܢ�;���!�ܿ�M�b:�84�F��	����N1e/��,�+c.���fII��<HX~��A�g���ʧ���fFJD��
(�#H��}?��'�ױ��>��jQ�����n��|��� OII�����M.踀lQ�q�b��h -��U��&[�3��5��((ue���H	F���ʁ�cʿÒYAg��ws�95A��!3v��یM���f����O�at�N����(�h\�l��Rq`O��U�a��z�T��:w��U��`'8�f�=#���!���WhK�k�籥f�rmgw��`�L ���� �L �ϘۧGlj�3W:�R;�CY�0ћ������ϓ�?=-)��JZ{�d���ωDc�@�N���v򎍉CP���P}�5���|�Ø�4�BSV��� B��LJ�E���G�w�{�P�������PGC��9|+�Y�}�9���ʗl,n�5����	��AyN��-�N��V�N���1� 	��A�I'�V'�m,��x�za�m@�r�1,̽�;Y�'xt3�ڠF�n/���\��$�7Y��jwF�[8,g4�� <Q�v�����O���P���V���zT&ъP4_.��M^���y�ԑw����]0⧰� p�DW�3�H����p�������Z�6_�e�'d���e�i�v�>�!'�<L����S@�#T��B�M�攫(��=S\�㆓�q�^���9�Cf-��č.dp���ǒ����NCNN&��jp�+m��C�`�O��b<�#�Y�fJ�t���n�iPՐ9�K��am@�B���K�Gx�4V�Ȅ��`������C�F��E?�=uv���"�E-��EE�#���w�j�n����பP�����ye�8w�o<��jV� =���N��G���?�h�C\(L�'�p���h��"!�P�m���mvg��|����A�^];:nxO�$q`|A6%�RI����t�ߏw�F�;��D��n��v}�ym5�p��U��9-�MpPaD1���`^�)�� �gz>��{�#���< ڮ������G4g���
=�,=B���&t�F�`/���ix��"���6���Enͩx&��)�S>����F��-��iKf�n���_8i�
����_��>�� ��JtqU��OӋ�R�y_��[ր�ղ(�H��X�����T�5�]K.�$l9�4��{z=h�AJ6pN7�+^�I���`�иt���R7�)����ѩ�񨊘���z�BJeV��8�%��9��qέy��.��IN��r�a�<�l�/�3&h=���l���EYq�4����Jׅ�-z���_a��K�Cঋ#\sÇ=m�8�1���^B�z!���P.>\%�fק�o���.)$�UO�Z[[���Ϙ�҂r/թ���F6v�|�� ���6�NG���������.�+��,x��Ȱ��¡�#���X؅�q�^�_S��in��ڑ:�F`?�U!~H�گe��kB�!�&����pu� �s�|D���F�.�s��06"��Wd-#B��D���s*F�.���~4K���14?A_K�Rfw����gh�{i���گID+<���	��X4kC��X/O�O(���U$|xZF�>VX��K�?���t$o�^�'�hz�xc(�K��A1�uT6.�>���GoB~:e�^ј�㨔�K���Lz��ǀM�1���Y#rʋ�s~QE�����q�_�l7p�á��{N���id�@�g]�CĞS^Ez@[J�DR0�U ��J��Uʐ}ǣ�B���`z�C*`wSԡ����l�