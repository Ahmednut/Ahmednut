XlxV64EB    1d20     9f0h�V湼�~��q��_�G�� ���R9��=a�T�� �s��S�������x��>�Yv�IY��(�IA Ǟ�Z_5��)oR@d��߁lV���N�0a����k:~�Ho�{��ּ�h�(�N1w̸vP/��wl�ش>W��a����`b����sM}�L��3�#������t.`��Y�kv��95С��#�o�\�8�x�z�P!"�Z;�s6�G�YS�5rF�� 0ÒF8�PV��䶒���ڪ��p7�ar*�*�sW��:Βit�IpY�i	j,<T�a"�G�
�A8�B���9��記�U4:���@�V�k|���F]*�XQ�I�-deK��^ٸ5�3[�tH��o9�D�f�{Ķ���W^fb�r�Qm�K����cS���
)v��d{��A����0w<b/���p���9��o��D��	9t���ʃd�^�Y),�:6��6�_a���eb���!�Kd:�-��.��m:ri�<�������Rb��:/������F��_��4����z΀ݰ��r�g9��,>)F	gjR�܆�a/�Ro� �=a ���*�#�O}n��=��D�0���x�Z2�H,L����0<SԸ=?��ҡ� ]]?ӻ[�a�7�<H��ZmI�}���?{?ǳv ɋ��,vd
� �1��T�Y�æY���u:��ꀭ�M}�'��D jE-$��VC�����L�������Ux@�2�?4@ ����	 ��!��^58��N�U�,��%
����<�n-x>�>v�C�9��Vښ+�n��A$p�yR�VY	���Z�~t�G���.�c�9Rd������K* U�tߗ�8 �(C;E��1�\�v��G��|�)Ucͭ�c���!�;�8(_SU�,'"\7���%æxyj�W9;����J?�ަ�^�Uc0���д7���&Q�Su��?U N(�?��7��B���}�Bbz�p��p��(�)cV`k*O_
�<��z~���c�K�w�����O���s�"r� :;.�z�&�����X�0�6`] >����m^��̊�lq����85����m)��2%��4�)N���6��[�d��n��^2F�U�6o��5&�oת�}��YP��w_�:E����A�����x���j�L�E�p	�1Tt_�s�0˸2Ki��B�:k��Vc�Q�?f�_8K����˧�$=�7t��K�:��-�6́�P��W%��m<��i��21�~
���tP���Q��D#%�$;�Oo�jd���b�k��Z�Iu�����T�T����s�� �X��>�d���ʏޫ]�Z ����Gi����9�Q����¦Y�+P.Z����&���Pi;{宀�Cn�)�"�j;cX\�^*����}O��rٲ����s��?�e�Z"x��"E�fN1��q!�T�i�jЅG��玢�!����&=r.9gO#v%�m��Z>��c�9��$��B`�=��;9��U��퀜���KcIR��5>�� ���Eʝ�?Dʱ��@�7 ��^��o�~�}B�SF���'{�b%M7yD_��9�|�T����E2���e:;�!�?���,r�gks��6����!��{	|����Q�x��r��?�.XO��kGK�&]���Fb�b-�0z��M��������������󗛥�O^���SI�؆k'M܁��!�p7��([��V`�\,�p��qm63jyF�"�}�<�ۛ������`s�߀�bg^+��=���tt�(�H4�Z<y[!+PQ]n|2�w}F�3!G��$x����_*�1f�����SԈ5SZ��'�ɽ5��㻱")���Lg%���u��ː��y�:�G��_��p��nH�T�Ls�)�.\i�&#��kv���]��]���뎭��l>�x]&�A�;1[�O*�DSq���S�h��s��ЦE�
�*�,-� �P[�_���f�lH� 3&�d1b��@�h5]�:��MR-��W�Y'�4_Pf�=m���V��ͅշB��Nc%e����,W��.��L\�4�#H�.x����zi�����ul#��:�xa�V��a�'}�yc�	ߘ�[8O	|������گ�|�	+�~Ut�[��쁏�UN���{��U��"��ã���&��7J������2��}U��|T?��X(�od��*ќUZ3l�f�bSU�h*l�����܇K5FEZw6�x#&�S(�ڝ&u ��I�0:��5���(�Q���z�Yof���ߍ�R�"[�;k��6W��{:��Y<�ΰ����ɞ���o�X��u������Kѩ���kh�&���(�q-o�m8���T��l�{��3d���]��r�T�8�컏en��P2����
��8c��wV!b���;���K�YRA'�.�6e��o[��%h��m9@����y��S�S�^��m|�פ��'�����I����e[7+��$