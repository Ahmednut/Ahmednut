XlxV64EB    1f6e     9d0D��� ��?t��~���+",&Pp6�p�i;!? �����n�u e�YIC`��܍�q�|�)����H���Ta�ќ��d�{޿��"ThV~ ��]�����`Ĺ�b�s�
c�R�1��d�K5r�k�>��&7�?>��/c���F��ڼ�Q�X���g��,o�Y {��	��1���Wb���~U��FD� xEmiᥖ'{�X�����V�xwj�����xĸ��?󪭶�Ȉ�o��yF��U���˹��|သm���l�C�<t��b������A������%-[�~i�����X��Q�*$���
Ĕ?��n�	2���Ž�ڟ����h9��=�-����c�,��<���T<)%d��ʂ�����oo��ð�@�&:m�a������ա=��(h�K"��|ݠT�|�s7�*Z�Ⓣ|�Pfh|F�$�]z׻c��G}�̤��V���G*�&KJ,$GӋ�wL���\阣��B�YID���(�`\�l1��_�s��F�����0i��y�+y]�)]w���8����fx�Dǟ�qDuz+�!��+�]C���6�5��3�(u1R;���kT}���Y��>5F���:
Ec��.O��$*)��8(Z�+��< {�~��9֧� צ���5�1ؚ���<
���Ӣ�����u9�,�7wcf�Pg�X�E���r��s[]��|F�O�b��w���NaZQ,,���O@���������Bx�%C�\����y��Quζ�ͱ��v�g^j�c�w '���w��s��<(;P�*8D�׽tcH���OU����:a�I>��	�CC����d�z-w��DU�4C��~͐�`w�++��	� �M��"��6� ZCa��+�r?���%M��^�N��>Zw�)�ູ��Lא!EMJ����&�_7���Ej�S��8�\^׈�>�������A;���Y��g���(-�]@-V�E�Wv)���W/d�;�7��%��O�4���N}HS.� �JW}��z�q�:z�Q��:���9���V1�<(h1~+���y�r�[���/��$�kH�0�8��w#�kF�7X?�W%֡��Zv���փY!0~>�1Mn=Ϻ�,�n����}L�&���{K-)K/�èj�I=��$S�������/�I�R��]�qj�wP�����H�K���Ǻ���UDX�/W��*�O�R��ts��q���Ĩmێw�Ć��lz���S�zW9LkFL�.v���n�,��d��5�؜5���2.
�H�Zhyy.�"��^/$�6�O�z���򇀋�:�j?�c�|�7B�	��4#Վ����t��:�{}�Fk�D]�v����	S@��lۗ.�x�:R�h�H�GH���יl�ܤ�s<'���xz�6Z���L�*y��sW�vc]��d �]�2���OQRAϚ�5Z�_�M��6"r�%iژ��Yw߇��)�;�X� ����N_ܮ��Xԟ���Rz� ��[A�HV����gU�=ԴK�����ٿw" S%1�V�}|����;����daN[p�l��_���j̰�t���[�C��J
|�ZF���KD"'pΐ�	� �@waru�c$DS���;>�xކߣ�ڙ����2�����4�=r�'>�hu���d�*� /	J�y������j����[��>Zf���z3_jL|���6�����(GdY��9��[�0�~ ��(��v��P4v�W� :z3D�&rm	^��~K�
�]�|�Cx�'%͜]�$�����W���v#��E!ڲ�\�9>cw�<t&UW��[Ms�wx�7���t0���nj�"	��#��~[�Ʃ��́�	Dq��*:\��ӯ��le�͏�9�3�4�*����[�s	��*�9��r��8�}��]��/X�@�m��� P{�C�#�r���G1��Ṋ�1�Gp��.b�O�N�)�����{�bAO����~��������y��;؉qL�]Ad�=����1�.v�:�ա#M�N�rd�˅��a~��-F��Q5��U�U��N	�/Ǻ��!J?��w]�؇�x��K���W$N��Į1
��~��ث���FmZ���M���H�����6��J��o��mni�i4j��n"��k���d����9l��o��i:��h-T�������2��:o*���p|;��Xz�8�)��������H5%;� �������$lK��f@*W	�y7����LX�=#?xm1w���"f̹ϲ���D�K���ة��%v�=t5��-)s�B#c��w�������<WY+H�1�Ym�G�i������Be��f�X2��iT���h���O��z�癘,C"����j�K�[�y�n݇$����[�j�٭+�_ I��ʶ��EtN��b[[8�K��Ox�s�