XlxV64EB    171d     870���i���2�F@�����"��r��n�.g���_�B��1D�eU��^��J���Q��ڶ
'�:�360��U����K��7m�������2�S�O��70�F+���\$�R�T�!�N�>����[,���{t#5i5��$�����M�{��o��˟���B�mE10����_ɹ�?�0c�u�5���7�����F �.�Sm���"v����0x��vJ�p�󏦺��Oύ�.�������16���yɨ�AFQ�K�]@z�:�V�$� �����{mߦU�w��� j ]C�ǈ��1���bȁ����ዿ�ҧ�?�#r��3C���#2H�
��]�(�v!c�I?��� ���c;�C���U����|�_�X=`s�8Q�d��g�	�bRH�_Ү8:�|glaw�z&��TN'vƊeG8� U�Ǻ -�����#�.�!�\���F:�	k ��toc�b6��b�
s�u Z�2���;�T�R��9��!��`!N�q�0�a�Z.\�$��ըܚ��n^��Ƴ��G��=v�Z��g��@qq�����2y��ڶ_!-aG��� �N.�>4l�6Z�a'���L4$�Q�qҍE�G�ͮ8r�h�L�ymD~%��j���NI0JMj�:�\��]��Z����M��1@�О�đ�� x(�6Z�8�C��5�i^:�P��qr��l��x��?������h�A����l<��ͥ�Ro��Tѡ���̂h6�H%�b�U�F>�s��ا!kXAzW����,^8��J!�<��J�a��0�D�\?Q#ΎNff��� 4�?��
co#�R��l��/�bN/O��뤹2�a���-A�?��r$���QH6�ɱ����#�1K7AJ�%���~J(y��iV��sjd��}��ՓT�0��k�2��L
֬2
H��qc��3��-�H�faF���i�n�3ơ�.LLY@��k] �B�k�]
�^{:j&�a�B߃ǟs����s�Q�� 6�x���y9bz����#��9P����#���yCd�Q��^��!7��p�05���51��s��P�w�w�He.�?�3;db��O�Oo�b��_Ͻ��o�"�����=��f�]�pgϧ7�wa)X�HM��.��Z��Neb�fλ�Ad#6��bI�v���	]+��ۊY9�ғ�T�l}�E�Bە_�ƶ��z/���C�7B�A��|	f�#u@Ծ0���k����1�ۨ���?�G��30u���e�-�W�1��:�wY�ȧo��7��j�`c-�+�I�,Wi�V�'�8��^H�ԣ�z����t��n%�Gà�� ɏVpF�pxYs`��;�rM+m"bMJ#��v/#<�trd��ؒs��1��2R�����y��üHw���(PeX�!}���r�%ϭ��n7�s�/� 96��WB��?�R���3~���C����aa��2H}bՇ@�b�ׅ����:��������O�CX�����ъ#+~���t-}s�ΡD������$����LN�շ���D��q�w��hg��a�� ^�D�N�P�����p�uḁ����U���`�%�%�?������{K�u/l�����n��c�ܔ������09�߳ڠ!����e������}]���D�V�$���$��#�sqZ����>D�&[ϻ\��6�[���Ļ���?�:��֯F��~�����|2����(c��5�/oc���#�1��~��J.kǈg(�k[U�8x`�1���m_ܞ�{yJ�S�/�*Iح;��:�/Pb��t�u�0�Ή��4H���˛\�����(X���ɀ�{���~��0��6?���t;��=|Ｉ�������5��œ.JU�P@��3�{��U�m�^zH]&�F����m3�:N��s��?a�|���'��WJ1U{�lm ��}��y	l���ؿB�?����0NH����H8?ܭpxl���e@�qRO���f�l��u���K�p���o�P
h�hM�*�w�i59k㝓�2��N��E��?~����9����de3t5����^�Tꄐ���a���a�e������<��t:B��l��p��