XlxV64EB    25b4     bc0\LT�U�V�M�@��ȵa���J��n�f��]g�_	7�u=��\1c>��1�2
Y��3�	���>�߁��%^��UCm$Է��چ��"V�Tb;L���X�;�4�/���$g̳%P�,�ZƍM���d�7|�-uSk���J��u���^L(dB���Uv����ｦ�i�C.mc�
��~\^	���z�{t����l�;X\/e�Ɏ�R>��8C�҃~v�	��eQr�󼊗�rt�
�wxڵ��\��u �M�������������o�Bu�!�����3�G��^��>���2i� �[ �l��][�P1l>nx�ϕr
QA]�ej1IY��EQ���I����؅�"NW�D�Yp�7^����R9��s���=�����T�&O��2��1��[��d��NG��-`5���@��t�zZɲ���)���2�IvO+
�O �1ԥ��R���nFӽ$����^�
�͸�_
=ibe��VI��x�?���Ol�]� �L{a�zf��nW�Ǟo���bB�{ ��aY�o����!g&�)��o�RLa)�ݺ6bl:���Z�4o��" �$h�@k�a�Nf��Ey9 ��ꃠ��}�.�����ܜ��Q�Q[a�|�N}v��1�Q��j
�I�fs�K�&���=�=�(6��C�fj�߆�d������u+̵��ՋZ��f�4U߈�:���+X}�����҄�c����1��p�S_ ��Sj��-��$�'������|�K�"�&:H�N �â
25e�&��eCc��@L��"��̋��-
� �D;���K�J�����R���Yփ���X*�A}OVM��6���v��#̍Vc�S��?q�#�{��z�6�j%����<?�Ap�h#�$	��(P�?�&j#Y�)���;��-��-E{�k��u�y��.�Q��m�3��@-T�,:�6���5�K^��y��?��w���� ��3)�ii�_�+";���mH���l�k���;p�;�A�qL�U�
�s�'�%��7��2�����+�]T�̣-�f.�wS�h*@��_�Ũ�'y�G���8�s�����
�^��f�wiTJ�a,�?�<��E��>����Q��������&e�q�aMq(7� IV�ir����������Z��U��ŧ�������FCrKT>B��VJmچ�2 �X��9v���e;!��<��re�mk"�]3|�kQ=��;�3�c��S�8������^��ٲ���}�}�r�7�.����V��	�	1ł�}����*��ʡ}�B6Y$�B=���!q�ϹJ0�Ro����V���V�ɨw0�!FtAO�18�<{�@��&Z)�LZƼC>ü&��l�2���%���n��hb��A�g���k��#k��x���j�-%�{�@[\�;�[���}#����\��éG��s��/�1"���k�Lx�|���A���w Oo��{��H�g�tCO�#9���d�n��lwERle/n�A��Q�*.�-����8jԩSj.����x1��jfli�Nu���v+֒��0~�?/x����vx���l��e��|����*&�/1���˧ {���l;u��ZS���2�R���&LA�,$�������S}o�9��^��H��$٬a��SY�+>�����7�xzǭ��R��UZk��d���^Wu*nj�<,C������3���y���b�;#Jd��N������q#���T�S�C	�\��df�}T\J{X_0<��c@Ӛ30�ΡU����B��R���w_~'�]f�����G�H����|	��(����zpz1T�`�wj�]E��t)�Wa,!𔠽�ē M�*"��͖���]�����V�?g���~�B��ekR�@c�|)�G�?�M븦��Sk�����g;E
q��A��0l����o�,��yn��|���k���cZG���j�u'��e��ȳ��8�$��3�H!�&����Kb��_�*v��ƍGj�t�ָ�����s�W�z��)Y�p���C�I�\������&|�XO'��ߴ�]�����A��_���)���C {�=_l ��m��(�pz! �4��m�II�%K��$5<����`3}���d¢HU�g1����o�\�����ʉ�/�������Z���V>�݈���\!���n���n�2�"����.�?+���Һ=�l�G�	���?�ҙ�6q�㗸m%�~��������=�F_jV6ڮ���C��Tq_�;X��@���n`�?�3ʝ|�i7d��NT�bP��a��es�>?�Sp04�Vw��|d�2�3pgK�����o�����̟`�o	�
�P6\��,H�xXfw��n=1r�tN&7=,�*��u�#p��mÇ�ُa���x����]j�˶aM(?�(�k�ڀ��LL��6>$tZB� ��f�MU��P�4����"�y��
|�����6�8$��o���y�f�lɥ�`s��ToFP���s�>��_𪵇ˢ��ڐc��kO�C����g����WR5�g�WTe��r��<��+E&r$�rץ��>�{"C�2��vl颛^\���[bQ$,G�n�V���y%φ�)��4�W��vQ�}L�ٲ����u�k\2X@2�vA�#Ч/�LZ�%Ž�R*�2;7a*)U��Ī���2�<�=)/y�h���q��W�w��pb�v��ճ�(<�͎r+s3���r�����v�>ȼ��"������bOn��bؖ��ճ��L݃�>&�*�$b����7m�T��!��*_���x"��y^<E�;SVὖc�é=E�����P�bAv�15��PZ�@UAD\�f�M�oU�&`�N[�[�ɺ�s� Ӌx�!��>:v>�)&+OX��fJ{	����#<�/��