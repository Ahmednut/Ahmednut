XlxV64EB    154a     7e0doe�� �ȓ&��{��e�T~���2���2ҏq��vVɹo�KY%��h�����#����= 7��l��v��ũSo���Mn�X/�
�!J���4����3����9�%4f��@�m��ț��a_պŉ|�l�����X��ٺ�E��e���Y
��/8,���3ҩ�Ẁ�[
S�e����i��d�%%�K��K��N�[z�y��ϰ<�7��#͕�	x����J���S�M'Fre��A��;����|*�-[�9_��7[)�L�D�%%�f�V}���<��Nfu?���?�q؋�3#��@9~<�E%R�j	��
�<��l��
�"�51@�=.�ti�Be7/M5��|B�ؤ�A[��=�Ś:|�=Wњ�t؁�s�%���+T�a���Y��+�>1�ɂ%�y0�ƾH��� 1��4�3*<эg �G���� ��gz�;7|���C�$�Qğ�n�Cf�a�Ty�o��Ї�B�$:���#8ym�ʻ�1@�l؂Kנ(����p���E&2��>T}�P�8N�� �1^}~Y)Ej�?��`�aC��*ٛ�%r3��c�-�KAeG���\i��p^��_���<`�e�WM�N�m�j�fik�
�/��3�('t�6G�Ov �-��Z�NBA��!�,�G��7�K�os��b��S�qȑӽw������y�m��'�3ҫ�zp)�tzۥӣ�ɥ����Q����z���uD䳓Fq�t��a�,�glF�K�V-�SU�{	)�(t�O�TZR>�B��c[	`ѳq�E7���*y���4R#�6+������b#2��+�3�/p?���gy�o���.B��t�_� ��$m�q�;ؑ�bp�t��U�����,h�[�����5����^⻖1�fw!L|5:��	[�0�d����6�����$2@�7��P-%k�� PjM�g�V4*3�wX����>X�m'�g6p��
@�m����Z^���ao��σW3��"��(*�����7,�ѳ��K�wo�/5>xZXje���IK�ɇ���^[Ɵ싍is�e�P�u(�A ��ԥt����h@��p�$�D�>��To�8��^~��U�����߃:����m�v�`��sI�t�T\Y�Ҝ	��[����>���/|����:QQi���]��x�M�ϯ�0U�tTwR>�zȽ��(��k�V�[w�w�b�gE�[G���֊�`"�� sX퇘�0��誜��~��G=��^kR��VΊ�O��/�,ݗ���y-ǆ��ػ�����q�˙�ϳ��1k�*�l��"\dq�۶H�c�2��r	�<��er�3\+3�ϝzwr�S���� ��\�;t���䞫�,�b�_�	7�l�M���WJ��AuB�g�N�O�v�7,wF&�W�}��*����je��z�7�FA�(��A���k@FAC��k7����M -3a�"Řc'.u�����-Ԁ.S1hmJ�;��B٢!&@�nt���7��	��>Q+]�k����S�d���1����"���"�������IL�3��4?�$\2y���B�f0U����x�_c�,@QY���"�)�£a�V�zc���=y��W�O��IA?4t�@՘_L���^� u)k҈e�b�����o���G���͉�EW�&/AD���������vʯ�P%X���遃>�w�K�c�y�+N��ɏ���p���>�t	�^�Sr��u[ӽX	�q�u�T�-�sY���E4���^��$�柢�[���V������ �y��?x\�~�XP�q
����{��mFkvt�`�"<�����J�Ap����lyB�����wH�����E�o�К�n�Q�ˢ�%Ͻ����O��eG�Y����D {<���eO�*�/p#(�¥�X��Tq�'Di���$�
1�Sz-V%�t�?��rv{8HPRh��_�ۗ4+���Z���yk��cC:��#_�