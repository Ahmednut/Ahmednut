XlxV64EB    6188    14a0ʊs�'�i�d�2�rZ�z���������?o�]���j�u>����0d� �}d�/flZ�?,�د��Їo�8�����=%�D������G��,[�/�q6
�����7`�/@�����z��b��ə��d�״N�|m��9U&�e�ovlBU�п�k��a������և�=
�7z��\5���������|�E�"݈�D��ή�u\$�QX�������:	�.e�[�Ǘ�+���rZ5î j+2��N��z�b�$����yaa���}��/�����?y�m�a�gD|��P�� ��$��t�����j��\a��ܯF~�fm�fD�j���Je[��0����?�)U>��w�f�W���{̙q3�I���Y>��%��\�n��9ԥa�;�%=3��fS1���/#�E�8��9Fe�8ߪ�D�V��n��XB�)�O4Ȍo�	@0X{�����Ӭ�V�Ԛr
a.{[ؗ�}��8j�n�C�M�]�9�d�4��Ɛb%��^��T��F�T�)ү���	��5ΰxAKjҞ��ZK?D1?G���piϛ
�[���:�cL�tI��Y�Y}G�0;f*��o<�=�:�x�K^� ˙u���'`����M����$p��d˘m��*�����n譠���V���uL+��O�6N�(t!��Bb�0�^Ԗ�A]�pR���f=���ό5g$�+�&,�����Rr����
�_��D���џ�-�!'��;y��%ٽ:��Zy^�7 ~\}O���¯dI���:v����?�!{���%��Z�QUU�U�gsܱB�qI�a������g�K*���Pb%Mv;A�*�q�g��wkd"�I��0�i���TV9���8�G=J��]֐u�@�yB0�L&�6��fR��^;� �4W�u�w����^�t0յ�`7�о���#�T�T���c-O������qya���q��fp{ ����}�ah�%��P������Ř�����J/ k�J������W���-k�X����2P:7-����:u�5p�;1 O���mJ3�����U�����-��%�5�FAb�^���waS���8İ����%,�YA�¿3#�:�!#+оC%�N�v)���T3�EE�)J�:��9S#?h�<_������:�S�������Y��ޅi�gAr����#9I4G,%�X]�A���v��Φ�8��=���g6�d���V�)X$@㬬�/#^"i���<��	�<�k+��X]�GF�n���y����?�U��&�=��4��7���oW�rIP���l0~���P�qx��׭A)�����ScK:V�8�z���z.R}M�料
�<��t"w�b���\�}&sp��;If��|p���-��XҒ�[��'m�[��t��d�s�Zs/�糰�).a�u��5)�r �_i&W���ZxR�x��[����u-�g]	�b�nyli�1u�ѓ]�7��Jω��|F+��|��fF������C����R<�=�/��n�M(wwͰ����G8[X�m�"CȠ��o�!�zH��t֠�͓4�\�x6J��i�����t�4S�v<j�%j5t�Q|u^��s*E��E@`-ӽ���+@�e�~m��S-Yg���%�_A��|�f&>�)(��(��0����� k�r��%#����V���͟;��FA�Aj�f��%�1��i��%L��T��45m�7��N�1�d>���Qe������1�0i7%4��k+J�Tp� �^X�n���^��'�W���]�Q��g�edV�w�P2���F}ܯiǧ����FZ�a�2��Q�d�l�m�Ɔ+��$+���(�6�p�K
h����i���6�l��m`�W��2U���Cm�Ǉ��<(|#^\V�B�`g�	�-�n9��`�}�<5�;E>���Jh�]�9����O����j$�J9�݄{Ϟ���Ro�Z^h�b�b0�HlԖJ�讙*.��C�5��r��b��aZﾮ�1���f���d�[z��8=N�o��\�:��J���a�`*{�ܞY��k}��YQ���V��A�{S�x��-X0�h����Ơ�;�,��B7΢ ���6����VF�!��[-�D�V��ra��Q��L�\ ��*�b$�oF��-�����7(�nv�]E���?�I�G$ru�P_�h�K���1����eEiHd)��4�`n���+�,��� Bc�}��Ƹv��z#r4id
�}���K������A� ��,��N1L���FT'gA��^��M�L��4��\}�Q_g�|�	ُ�e`��Ǆ�
s'$ �й�Y{jw2�-,@��gL������i�Bj��?�r��oė*�T��/6Na�(�i9[���*�lm�TI*������sѸf��,`�*�D71�v�ӓ\>ik�J����VDay�J�"I��5���$���P!�#Ö
��^#y}*��7�E�4�V�����R����0i�[K����:-����v4 <��>B�{��L���	���$H�����R^"�:N�'���^��S��z�v�����N��hw����[��,%\�K��i����9D
R��}�)�l!�y�π�6`��A�����K?:����n��$�@���ʥ^�]�����~h4�����a=r_�
���Wo<�]��2<u�[+����e�yUJF��S��*?^�]�@Z�ޛ�pW���5c��3X�;�:��~ٶ�ws�w�U;۶'�3���1 �a�C�f����^)a���(�^&
�t6��"���T B���Wq�]���vs-5'���-�0ը��h*�/�(�mD��G�c�E�ן켍w�ܬKƺ^d*��$�I��W�}s���"�\�>|���\i�!B7�F�?�PE?ߙZ�vgϗ	��m�����K�0y�����g����%o�����q�J�Ⴉ��q}�8v��f(/zG��7�W��QwqE����v	���N��#|����O)�|LH��0�ʁ)�y�b���[�U�P�P2<H��5�FL��+�uOyhU_�
 �᝙}�%s�C�<�D/$��񷡔
j��lw�[�������H"w�
�B?�� ?����}��?a��<�\JO9�9�< 8�UGU����"w���Q6�ZƐ�w{!�u&A�gӻ�z�o.J<%F+�囌��C�p9�K�:?��^tέ\�K���^#T���w��9{�����Ԁ	Y�)9UĆ m�$��^��H�+O�)d�0��	y�_��q^j�R�C�۽�	��7>?و�ue�.�:}���h��]BDЯQ�YU;Eh?"� ?�Mf �R_���J�\4Q�V����^�����^ �+d���
-ih�ό��bp��=h�B3�����c�z? �v�:�
�h��@�AM�n���C����ِ��s# C: �?qU�8`�\|�֩֫���n,��b�EB�]�E��Wc�	@�#�QxA*^=H��� 쟴V[<�θ]y��)hD+d�5������bmP�b*�$8��^���U����P�drۍ����1('�r���D⥴.I��U��C�������j0尠��Ll����8����ٟ��$�5�R�b�� k\6��m�] v��$$�@������p�̕i6�LE(t;{�Ӣr{`҉�i��-�ն���B�[r��Ƶ�f� ws~pR�kF)�<� �7�X�F�Ϩ�}��@Y�v�ϑ��*�=g�}U�zԓ��ɕ����z��9+��_���{=�B�1��D0�	��_�[	.��w��Y�Y�~Z,�J��DV��Q���`��/�%�zA��v4���2�!��Fײ=%`'�+6��`J����5���5ƒ0h�CW�&�iT$�S�ޔ=�`���D>�
��6���|�r-���	T{��7qS��:͈�\v�L��[
j�X0˷�Q�a��vi �S>J�h��
N�1��<�T�2�ٿ��_�*�t�o#�8�C��YY��`4��4`b�����O��u�=��	`����9T�P~�>�)�����ˢcL�$�D�?l�ҳvjE����N~���C CH�_���j�O{a�dq�13��v�S�4P'���dKA|w&#�*5�$Ҡ������h�~&X�k4�/y\�e�ᐼpՇI�k�Q��_�VV�/����_G����Pț������eY�\6S��j*R�U�И�Q����7��;߃�8y�����فFQ.3H����QPju�eO~E�(ux��k��Ur3�e�ޙG��.��\�������Z�o�{Kz]މL�?����˥��
�Bv��._�����i�*��`��)y�����\-� %�g�D��"��YJY���
��)�a�s���B��j7ш�U$�i!ҁ@��7�d�d�ұA�B,x-������)^rU��u\lC��M��.3�G&�"e`g�U����,H��o�cK��'����P�˵D_�a% Y9�?�{��ޒ�Ɨ�'&J4����?����#��z��e)�w���آ�8�F�"�B�������r]Zw[#�m詂%��~�>rR���M.��&l�z����R�qg KGw�ª8uJ7��_�$��M=�$*ȃ�kw��Xs�o���_��jIw���G�	��u9%~��nYI��b�X�������J`u���[�:X�H�Ke����k�C�Bg�{�w���d��.%0o��w�yi�a��7$O*r��9�@B����"�'�]4�/5J�K���9l(����M�,�J=Q�!SHa��ڧ�����L)B.2*��\�;7�		�����f�x<U�2��� �I�CD�@;D��M�E]���[R��J����XS�����C:*y������1v�� �)�\+������ރ�3N7�B���z�.?ل��>5*u�8\��#Խ%��(]�yt���_�D"I-� ʽ����W�(0�N�p��6�u�����Yxl(AZ��J8�J���ߖP��,m�$� �%��>� /�sj�X�ث �0������|]4�~"�nܠy�F��A��O,VKh�cт��{"Ѯ�",y�
�1��h��Ɔ(�/��
\b�g�u