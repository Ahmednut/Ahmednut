XlxV64EB    3eee     eb0`������;ti�/�AB�$A�#3�HV.n#k�c}b�O@�X}Z��]>ܣ�9��#��0�u�&
D��O��ig0���5�h1���ň��>�H�V��l�S�0�]��)�u��=_��s�N���gZ�R�J�&F;p�����O�h��� �\�J�/dQ��L�T<^���,~�%$=4�ZFhtV�R�G��G~�r;�^��8�ў�-\ �jv�Ny��\�����w/]�^���
z c�%  ��ͩuz�xS?4ː�>-��t� ��?7uYspP�Y�f��Ν�g��V�'�6����<�}���(�u��6�:hIϓQ�N��8^�[1��UGw=
�>��%�++4l>m,Zϳ��j��'��S Yy�G�(V��.��m�� � �a�-,I½��.��̒`q9�p�@	H	/��~�/0E�Td���ϴ�*k��e[�_h��0r'��^���f�A3�:K�G�
X-��C^.�W���Z�^|0L�Wm�BK��2����e�ӗ�592�q�K�!J��>i�Nٔ���`|8?RJ%�q�����`���ޅSdl���迗֎��h�t��{
�n��+�}Xe"�\���i�}�y�|Q5��:8&M\*���>Ma~��]Ǧf�u��`�\�;S7|Ŵ;p� ���[%�ۗ"�(8B�H_�w��;=�d]`5Y��?B�I���^9��	x���J�S�T#����	�񍼲�F73Ai��!:J�,ӭ�3P�W4p�z3�du}P��
x� �g/��(���$��r��y���} �@$�%JҖ`�N����˾L)�v�d���H���)��0��}ֿ0��Ƭ�d�%�bNF�LkvX���3"QI�Q�条�zAbA��7;�/���� �ܾΞ[�u�m�v>�/���#e�6�Ɔ���s��X����Ǹ
�f��.�`��*���S�(v/f�"�Uh�������~;��l�3x�;h�W<$��h��}뒌�w�I�����R)�»]I�'pĒ���8К��膙Ը\ڦ<�٦���3o_@!vH�Ѕ�ס�Ew�׭`ƞ��$�]]��j���E�:,O�'i�g�_��^ !��w+x����6�L#׏�9sq�i�_���9�J�U���CkM��`o�ϒd�����}���5�#�b����m�����U�0z؇�������m&���듖R�۷i��@�~L�|�N !JY���c�
WؐV�050���Ȋba�rm����н��ޚ�
��2_w����k/���Ha��<[��R�R�|p���2a��wTk���A�kev���ԍ%���E<J�=V]l	uI�=�"4�}�Q�I�k�ʼUۺ7�Tpmq��`^a��M���=̢��Z�*�P�c��Q-�&���7�	��A������W�x*)wQ��v+�|bm�葎�F��c
���&DI���p�g�0�Ecdv�_�-�s6��aP �/�p�| yǈ;(:��=
 GӐ�}�7�y?��WK�6��SE%>Wb)�f6�.�C ���3.����r H=�Q�f�%�>���Q�&����F�R2%����2�a�����u�kc�ώh~~s�ֳ�A��wX#�sX;��~����:��<�m#�͝H
,�.s��`S��k[�@�e�� B�ү�H�U�o���ȍ���E�)nZ��-~��8��� �-WpU Y��4�O�A���� �#�����:�a��`�&���:����MQ�<Ff����6l���W�<71̬{&2B��$��+jǠ\o(�J��@q�R�ػ\A�B�����qYHM��sK9�"�f��_HaʝK-��	�K'���w�
���O�<��ԟ�%XqQ][�Q�!!�cc�7Nr�q����0����0��@�DB�������r%��B:����d`�\�4?��=pTPG��jo͵X_�d1S�.d����T1v$������R����w;�A� ������$��� �e��p�G�� �6�N�%h�cJ�?��u����ޮAv �]}�����3�><���#���Ͽ$tY��è�KBVve@L�KpN�٠�Ɩ3�0U�pi�`�{��ޟ���N�L6�I�U��Y�����Lb3�o���D�����t]A	b�L^�]2E�9;6,�G��FؐO�6+��ߌ�N�aie!H�mzҀ>�#�$q�*��5���b�qZ����$l��_�e;r҈�f��C8`��q�s3�"b�.�iK�J-&`vP�R"ot8�!�
�-z2����(ڣ1�W�SR�u��i��7�����L��|�7#�3w�h���4����Ɍ��[k�E�\���+o���5}I���F��=������Q�!�r����Ŋ9(����d`��U��U# �K,O���Ti��'
 {m�%���8�����yt?��ujxԢi�N%$"#�D��C|x��-С<��p��i2��hZʳ���2@T��I*�Ċ6�j�9�6�Q��Hc���F��W(#H���QD��H�Qm��W�n�
ùtQu�Jk�e3��a�b�_�ׇ�v�,Jǣ��r���B�m/N9:~j��m�r�6<�C_���.���͌���[��h𦧥��2��,V3�J���4�ƝA�?&�K�
��[��md�F�̊>�u���2b���Ƚq��XH����So�ߔ��d_?��k���H+ �
i0��i�4.�x$"���g�҇r��7�l��.�"gL&$w7��8�-�3eX��F%�dv;?�z@I�[#�_"�st�9����d���y\󌡉�v�˭�|����n$�]�O�+5�ƌ�V������Q$�Z�Ȭ����yk�X�!|s�� �7�Z�����4����ߙ+�|�@��k�t��!sX��Ӷ�&��3a�҄P�~�1
о����f���b��X����N��f��C���ro(��^�;:�����D���.8�Iʼc�̅�$e����vl�;��qA0�BC�d9�cKvh�8�|=;���G䖕�H.�+�F�3�X�v6��~�s��	�fm��D��1���^�r�ܐ.� ��Pqۇd�w���|���ぜ��R���<�h�x43��g9e�Ff�1xe�$4���$_��BO��dGUt��^H�fƬ�u�~�r�cCS��"��&�G�V^��u�h�:8��wNٔ��	��t�C���4l�>�8���b��Z��ɟ�s�(���0�)pQb�wH���b��2�-F���5��E���l���N���F��sY��m.j�48gz�>���WQ
����4�����\  �¥����I��2t�Pe98`��)���VZ�jsr��(F�5f��UP�5S�;�"�HN5������9}6�H�yǐX�ﲐ8.^ؙle���hM�!���ԐЀԻ���'<C�g���[�Qc�f���Y������=6��|w�%�Ղ�c����C�ϲ��Y��9��*�����8���s�,�c�B�v��$\��ϔa�6'5��N�@;�S�U�&8$�~Sꆡ*(+�����RX��V��H�SyX�<��!+�P��g;�*��g���&;yOP�DLNKۺ�}C��|�w,����/׫e����������t����|�aA�6�>%