XlxV64EB    19b0     9b0�)����(�~`�� ���c�Ƣ����T����Ʃ���o-�.�&0���*ﷇ���7"r�Z�J�(&�(���wQ=�d|��5sΟ�y�.�5��ˤs��m����W;�ќ�Q�^dkTJ3��mBD��/2�;�b3�Z����B��؅�zJp5t��WlĎ&��G�;���`���JX:�[�Q��iĚ򔹈7�c�҄1�`�
�_���+��n �ϋ�/�l��a�z�f7 ��5��"?.x+\M�]-2.�^�%ځ�q�M��� +�I����S�v��O�:f�ɜ��R J�f1����f8�R�*��lq��Z�A�H��b�B�R�ډs�Y�G$9E+!�>��;m��6#V=`G%��� ��p�؞�G����Q���K�PY}�(��c�7�\�;�C9����K��L�C�I.Yݾ�V�42�xv]^`;��3x.2X�b�O�(l�g���YwC��k�EJ�#�hl�.�~�n}���=x%��NK�m��.O�f�)-sz�Hh�[�>*n��ߑ�Vi��(u�g��Jݞ}��:��(��o>6Ƹ�����9��B���O�_���օl��%�[�^ŷs�����/w"]ۭf�E��Dc���Z����1�Fl+��q����f��+�����l�Q����'��0�%ik|[F�abL���-G�°��b�;�ZEz] �� �nC,�R�Vk���N�a�4��Z�E�A@��&��}5f0ژ�l4\~�%�@s�m
���X�F����e:��b��,@z�i��t��B"gk��z��L���@��x��צZ��i�2�㑙�NL��o����D �!)K�����An�f�|���j@�����)�!��MOi@��iU5Ǡ��s�aʃ���K鏃B�V��Q���,&���L4+fi��"A��O���?���V��(2���0vkn!��[=2��Aר�wTX��#����33�$���W%~�}V�a�'������]S��y=�5��������;}/����w� OQDڙr�),�5��?s>5��	qe�6�p��m��9?8�2�8@Hӈrp+�)���ز��R���&�ߡ+:(�[�xi{.�94�Y��يJr�ͥ'��v}	�ݖd�N,eӷ�ѴU��	�_���
\�A������zL%��&�A:#lW�oN�f�2�,+�x�XC�t��{C�H���ŷ0j&����&�㼹�
J�Y?��֪#�;t���� ,kk4����Wh�Ar(���Yߣ�"�V b�D�yH7�`
λ���^1hL5%+�3Ԯ�D�?eD�����z����m/������Z56O�5����D��=��n���
��l�J����ʻ�6=����-�`���d��n�ij�/39/��{P"t�)��7{��uU���0�7�^ר���b=�:J��Mkz�՗�_M��cRgG��s�y�=P��e�����DEz�ŀ��K�{u�Ҍn=E��Vv��]������ء�t(B�#P�]v
���2��p�OPKD7�V�V�湃��K|H�)A#c��������cL��)&y�+�z"ġ�
s/H�0{�U�R����}�6���������H�vA�պ��v�nH	��y�o, R"!W�ٶk��ŵ����d��� �
��|d�á+�^�hR���!���N�s@�P�YlJ������t��kw���#�~�B��б�d���Q%H/���fd@��g��"ؠ���P�KS��+��y�9�v5)�W+=�V�c_��� v) ʼ�i%�m�Mڙ�o��)��	
j֠A���J�C�0����8�S��΄��/���}�E7lxo�VD)H�HL���A��r�d~�����:�e���'�(c�՜z�H��As�n�͝,(W*�xqt�?)}R�J�z�5��	Z>��&���û �~g�������˭��x�8�A�v�U��47����	��NyCbQ,� �ڨ����o7=�Y�|F�ypT�K�լz�i>`���>���d��Z���µ:P�h�lY`�m	�����m~����V@�H!)s����R�kP�Ǽ��CZr7�`J^7`��а��(ˍ$�I%|��4��.�(��z��"�n�<yb���f���������-�7'�Av����W1�8�����}�@R��0 �9�/q3��L��
4�K��|�ś���̝a%V��n#�=4bW-a=�c������L����J�{�b3����X-&޼��n=lA���W��t7^�]�R�u0�AÓ�9����#��m������wW�<�� �T��Y���S����YS�/T�ċ�'2}E�[�%4��m�,۟��|�=�4}Ǎ{$~�}����Qe���{��oP����V��Bp��>&����fo nh'Zn�i�PP�C��b