XlxV64EB    fa00    2d40nЙ�#Ӳ
��K�E�DV�&��U@��Z�+Qz���-BKUx�����]��B%`5)��1v�s�k]�;	�'\6�����):����u/z	qV_Ɵ^�#|N>ٿ�&Y�U�wW0�H�{�}�e~LM�1���}Au܀��ր��T����f����42ay���	�$Q~*�k|#ϥ�F���S�|R�d}����Ҳ%yԭ��$F[�T���5���!+�����@HV˸��"Ir��D9�ߪ>�^�]?
#�q3P�5�JA�*��}���+i�Mh��%���_�"��_��9Ub��� 4M>?h�>Ӆz��	F�A�MuQo%�HQ�69��>��y���j]��X��$�Lv�=��e/L��il~շ1o��-���u�a�0<]��et���}*�g�:X���ݏ?����B���T2C��V�\������O���V�(�`=\�I����zDzL�M�����KhDhϩ��Z1z�N�Y]\����D�M�`��^a3Y�ʬ�˂�2UW��
������5߰���F��E�1$|�%�b+G��xk�g����ڲ~�b��_���(�m��	�鿦;��\��};�0q��$W�"�������X��w�N7��E;�Ǔ�*`�(�A��5�Nds&�F������)R����7N���@��M?��q���?�9.:D��^�c.C�hI'���w�;�a<�_@����G��'w]W��v'��hH�^������r�2�r�
'R�dU���,�9�t<�)���>�O�i�l�<�Q�t
���l�Qz�F�^��b ����
<��]�|lP�P*��g��	���0[te�ӧx|�����ʏR�m��a�7o�d���\�yr�]�|��Tͯ��g|�%���u��B ���Ӗ�7Ȩ	����4�y�i]���L���e&��(*�l�p�bֽ�;�q�/S~���#��o�UVK�eӍS&���vpKȸ4깄�kc�?�Q�,��k����A�����M�3D'v+ ��Ad�C��Dy����dlz����Z�Nl�s���R06�n*9�*��	V{*s���]?��_�H��K�N�(1���"�����V5Of�ojUKPM3eTO��c��O�d�]�5m��;�N=���bנ��=��iiض���(�nK��N�F���!A��>v�Zv+w�l̅fmuF^�۾���J�U�C�8W�I���nk8p����yZ@Z�ˮ��#�Vq/ݫ�g�^�	qv��<I��}�q�!���M�ϯ�5���5�TB�gU���������60���>dgm�+�,U�ߢ {������b_f�U?�D�t�%��`��fü���|h��':��u-}����kG��B8�}Lf'�y�}(cEvL��F_���"y�"���ݲoyy�X���#c�i.��-�[��/o�.��3"�9�Ūi,Oa��3�J�N��-�k��r�&4q��O���f�:#�2HG�2�S�V��s9��Ϗp_���y��%����τ�O�9_�^�%�G�|+���Ԅ�Dl"�"=�u?��;��K�7�� Y�ތ�<;�@��'��dcM�s��=L���
J鑯�&n/|�)j1x��{�8�r[yS��n�h����O5��;�s4 1�yuB.2ZP�k��3B!�F������qo�٢���� w��W�*<��9a��شJŔgx`���ܜ[�Ԛ�r��M1�\p��Dv^�qp�ew���jp��;ރd�.
�����9��_ ���BHsR��� � 4�+�Nu���6p:h���G��N��Qթo�;�O���n���b+�.����p�^`���\�@
���8t�&�Ȍ���=�K���
�.B�+Lt�y���oX>n���|C&�m�4{��2�W�n�q S����Vl� 
�q1��~
r��4C&3"_g3�:�#,vB̮
��`z��{a��o��zt��;$���y��	��t�E�D�C33�wA�}�!��x�*�c-H���P,~��?�Ek�C�]������EÌ������n�<�	!��y5�./�3c\u��&�����!�_�|q��iǆB��܅��;O��+@ݑp�ֹA��@Si�A���|Q�c��$aL1�,a����*_���b{��w��0��}���\��=��,!��#Z��r�@�.��@����̧������]~��j�IA��܌�����������Gw^�]��k�z��,`Ǟ�b�s�]�������I��3�M�zA{9p���V>�2�/���q,���D�q3���ۿt�(3�%�փf5}�l3D�	�N��2��O*E+9��H�8�v ! ��1Y���o��w��]
�T�K�Y���5S�D��<&�l˳��;&BH�|"�{^/Cmy�*�e�G�����uf,� h�P*Np�2ŷw{G`d�ݥ2��^��m����˄����읆ܜO��v[���*rʞ�`lI�izh�ƻѣs��v	��=g{͉��9$��Xc/� ��V�wg
���(=��;kk3�j�bL�I����İ��/Xk6J��Q�ZF�ؘ�	^_��Z?6�x�A֒�����'�"H�V���p�n��.�t+��$\����'3����a��dG�M���.�$O�n��? �9�l;J�m�`i�3��L�\m�8�ݭQ
�Q�F���Ƀl�v4nXXy> w?N��cv�䡑F���t�5{���(�2�Ǣ��������_�p�$�r��
�LX�o����&!>
��s��A�Ɛ{�����X65��U�e"a�
�c/VG��"�/.��-^6;,c��!w��|n*�*�b|De��L����vS������M$5"bV�!a�_>��p��q����K��� ~�d7!�S�,����P�cUczN��r	�z9���t�x�%��ѠX{�{�����ѩv��ݟ��É���|_v��m�Rk������U���;�[�#5�nb��on�1pd�)��:�g��	Vܦ��`b�g�%a��HP55�E!���k)�xm�G��t!VH�f��H&-Pre���bX ���`Q�*Ga%=�F ���i�B.�]M&T������y�:C~
b��\[�Y ��C�+��į���.��F v��+�5��Z�;50d��@�Z�@������X��6����qha�18�����#�pK��ؖu?����Q^�Myl�bAB&��t���^o��Y��5�Jq��W����ڡv81����[�B���φ=�b��_:5#����-�(ל���߹M�3���4Rx\g��y��U|YP��sYŭv��D.�w*���,]���)�����=>�I`o>�a`�I׷��f����^�.�iÙ�YU��F~�}E{Ҩ.G�k1/_��o�����9o�������,�.H:�
h6�6���R���.��H�<V�g"L7϶Q�n-��J�#��MWӐ�w߀u2)�<���T
Uku:KA~ sm$�	»P"P k�1W&�F��"�N/S��ߤ�orfJ��K���x(��f��k���db��J&����cf�],'=?�(-R��ɾ!K�O�9=���+{��ki]��YV0�؟�T-k�3��p�ZP���m�\}���ͦ��2��\����
Xv�/zrj�o��祴�uN�|4Z��%	��a|(�C:���W������Y�����|�Ot39v�����:��;��?��FU�o����K'	�l�#F��HU|�a_�1z��_}�d9�m��#�F����B&Ta���:��9�#^�ș#p���k�Jn���)J��5sh]ȸ�y��2/��I7���g\=��'��.���a�*<�ӣ_���j������0χ_�J�OkJiٵ�X'�W$C�1������\	�w�����1z��5z��{�
JV���lշ�+���&�}�2E}��ɥ�q<g4�x�s��.F:�\CK�Y�@y��+�qX�Y���	mN����~Y6U?�\���8K�ۗ?8@��C��u~�3��b�mf��J)[?��_�$��g]:_���SꝪ��-��X/������U��N�֏U�0q!�)��hb4��HI(J�y�ٝ��HW��`p[JC�ř�»!Y�#Nv/21款
'��X��҉Oe�p�V���� o�
��89�|e�̔xk9��8`z�}=3�q�x�IÀ��T�J��6o�S$[��/�� 0��m�/4#t!�4�G����߼�`�C�`ifZ�#;	&�&��=ρ��1'e�F�ᚵͅ����B�g��6z;.[� ޮ�'>���d���+�`h��$����c�[ٍFa����S��rh��o���R�JdS�օ�qn�� p����դ�NmXր%v(��Uf>�,@�G�����H86r.l��#)����y;�4����k���S� ���4��>K�q�
�������±�/4y�Uj���< �-�&и�n��|͒9�ǌ��W�/��lʌ��]����$5��9��3��M	�Χ��ÅB��u&��E����8�^m7X���������Q�u�D�΂�t�ް![�E����b6�x�qdîE2�V>0��HOX�=p��5;w0yW\4��������7���?s`�T�����ʻ-?��M]���Ⳕ粣��1��$��@�)'N]^<����2�E�mh�l\W՟�K����yv����Ě�ܢ6{3��+'H�yS}.���4v^���僸���B���}$];����Ǔ_����I��ٓk���nP�(��4��៣w�F��i�8%��^���B_����#�k�PX �4!�u�H�Qz�6�Y��|�R�)c3l��z�21����	Q
�4��U_�L� ��#�Ή��R��u5ht533K���@��W�z���]���uR���$b��PՔx�4k�@��Qz=x�kG���=�����6��(��t���@�[,q[����o�J3C͋D;��+�W�]L���D���@x<`ߧ �@3Ga���L��@�+���������+��p6�ES���ˡ��F!�X�e6�if�����@}\k������i�rM&)�#����`�szGH����v'U��⬹��><PdjT�{@��y(ގ�ˬE����U�z٪1``lQ��nӉaH��0������d?g�w�K�L�A]�N�:!qj�����I�"�4��KGљ�I�
F��]���㒩�4Z��������.-~���v�,��7j'
EG�{�P|���^F�qL�>��){ھ�J�<����c%J<�i�ynl��[m�Z\���j���i6M���15�TB�׊�	�Ya���S6�~�Aޠd>���Vp�j|��rYZ~َ��v�H�O��W~���#�(�J�q�c�i�����d��i����p��ӭ=���h1�:s�ރ�臐0��x��U9�O�E�[�??���.��\_FEPΏ|�
=����
Y��!t�Gq'�`�MMS)�"�2i}0��0]�X\5��U�q=֔�`��������a{E���N
�+Di��81�E ����!3�`�m3Σk���z�7�}i=�:�+�JB�)��;o&S��Z��4��Q���5��pA��-H�0^'�,���.�2��yxj��tg�4W*����4��1��vyO;�\���8�ۙ\�+'
�����Ӳ�l1੕3��x��c]p�-gs0�2nbd6����:�����b�)���Y1 � ��f>ClR�;��Y�ۺd1f8
�����6�h��k��FZ	[t���T�y�d�
���=>x!)�YCWS-��~Y��.��N�$�
~�c��`���!��~�[6]��Sw8�fmM�1���J<�Ϣf��Q���A�p��x��96�=��K`���B�j�d;��Jj���x�D_	��g���Y����.�1�Y`��ס=gG����\�}��$H�:*�>{�(n��cm���51Vl�h=E8Hf�WQ˷�j��+$/���� �.t ��(��4V��Ml�����E}Vza.�L��l����F�ۻ�/Ğl�I�K��ǃl�ˮ"��b�i�9ǔ��.��D��1�JE��c�׎�h)c�<�w(v؋a'@wH�������_q���X"v3N`+7��L�f���ks\��.g�@"-|��T�JHDPN�bF���,���O��,�{�3�T�����}�'��%T	����^RLV-% K^	cM���x�/"xy)h��� 煐� ��4��l��]R�j�z����\cOU�l� ���`���wY�I;� =[���������)�5�5PF�%�-����;�B�iQ������ms��t([}�]n�~�;�!�bmO�tH5�����x9�a�#r�������8���(��Y�j����֕�Ӗh��>�pGEv�k�XA����H��Vm�b�^��&��������CW�G��<�x����գIMKr�j�IXět^0o��O�7���Ҁӳ�9I���C�](���)�8�u�Y��/�z���:#�jآ����a�[�mVI�� o.�В�E��(��ͫ1��ʥ�#��%4��n�Il|���k:�p�4�"�Ju�%NrG3מe���c�C�����{2�Ko��#��j��T/�Ek�k����NY��60����؈s��V�&p�$���{�����%˿�����rN��c�����s�f%l	e�>���t K,
CvS��K	04-w�勲U�,���}w4^]ZY��␣3��%�:�(��ki�C���(P�Mp���A7I^/�m�>��S�^f��&W�c�Ŝ3��W����J�x�+"B���mE@��v�T&��׶����$ڬ�~���݌�i��.��mF� LH�C��x9T�cw4��lƃ�G�����5S:d��~�:�{l�qMilY��HS����*�>�`�N�q�q��[iI���@�L��Ҟ�	�X�1����2����[#ݳ�N�67�ݩqk$"C�Y��2�ù���^% pU8C��S��<��(4�]l��2�wqF�����
o2�j���������e0V.Nf#��Y��rAJ�)��	��՚;#� ٳ~���v�AH�r��j�*���{���Bk&K)�h�o�)or����-��i�oE�q���1z�f*c��tڲ+���xZ����kGΜ���' t�iG��c߃��gz+^��I7�W٥��%����-�V�a�m%����T���Ǝy���&
����ȴs���7 t�}�q9�=�&jh��2Ƈ|�n��b��j1_'���f=ݺ��t��#K�8^�I]Wτ�,UİU�X���X/�O��d%�L��,�]��7V�G�\����ĸ
D
�헆t=HN�6�D�����7Ȁ��{Q�w"��7JS� �9��^!bާ?��>��ƌ�>x�>���."� L8F �R'v�*�R�貛��HY
"t�׬M
�&��� s#�IK�"k����M�;B�Jx��l�1ܲI��� �ݳ� �ȃ���Wb9g��d ]�x�Zb��vh4���*��p���1g�	�� <������b����m�L2M�g�JP��52�G6(1��%�|S����M��; �Q�P��Q�����B��i;v4�-
Y�-�W&�|��J���!��U�$-v��P���5, �ގ��Љ�N���m�;��b�W�v���������\wK���L�|����6�ҹ�=�-L��u{n��>���/4��?�u!�-���B�H��F��e%�� ��w�Қ�Z#S;9���C��N� �Ƌ���(G3J-��u�+"�,��c(X��#x�7�(1�z��lBʦh|��!�%�U���v�n�ⷦl�0Z$V*�j�T�Z7/L�f�R+;�����iF�CR��ρ�6�BU����yp���D�$MӨ\I���ģi��>���ku�Xoj��z�Fh�:OM�R"͍��09Mi�ڭ��D�	��/��3dz�a|2���3HOe�a<�-U�Dx���xݢ�,'�ԩ��}���וD~�E��L�	�D�2n�ZVc�IJ��r���Buk B0f(�ߖ�T2���K���W�MK"�Y��"�-����F�����<�Dٶ���)Xn�g�Ƥ�����U�UVHT�d6��*�Ih����7�3�z��Lh� ����^d<���4�ã��I)ھ�]W=
�^�T��S�#;:���Z��)�	�B�Y�E�`���l��4Pd��:���'EG����/�����L�����JD�\���,��5fZū]�W-�t(v��*4�fg@xc�I����S!*�Y�5��'��p>J�w�F����35��7���%K��)��yU�˗�F��|L�=L�Nm�(������JK�/�p �#B tk�4MpWh�d��x���G�=��^uv�Vm�����a�w�3����iu�� ʌI��ɻ�-���
m���-Y��&�fp�"\$��'�rR�%}�`�����9 ҂�5�L�T󈃙���TTv��5�вhxJV�Ca�[G�%*�jti���u�4�.�>b�vi��������#�Ȱ�Y1!�lO�sc�+�r������3}��	L��Lk��ƆbiZ�E�Q���}/�y�Z4Pߒ?��$�l�8�ن(C�7mD��Q�.�1Fd;��{I� N�q�z{`VA�f{d�>y��(	n��Uܧ^G����=�P.R3�h��?�i���Ix:*��!����i�N|k�QkBoM��Ek��S��3F�¨^@=qÉ��<���@qT⌹�+W�!�^^T�����1�`F���;W��g��7�ʿ�ZG�J#�-�(��������|��7+�W��<�H@���H���<�]�AA4LsP<̖>�v��iq+^[����d�؟g����T'�Vcr��H���D�`�q�fFH����,(��Ὡl��H�X����&��T$p~�h*��'��ջ�&�Q��佷��1� ����K\�U15��m���yƏ1��<ۛ���OJ/�u���r"}�)�ma�M�b2/�	[��ob�����d3�/|(��򏑃�n�~�ux>l{?b8�ӗ5���#�( �͡{ڦwj軾A�9o�r��KT�[u�.��?6�&�e5?��,���9�.!�T*�Lpg��йc���PҞ���G+#��Z��mt�Ӟ� �a�,�c_��b����l�q䖄Ȋ7)^���>�悻���0z*I�3N~R�#zS�V'�K�U>ٖHٯ�Y$�B35eL7VI���0��T�8s�Ϫ��=�5�=<�]q�з��W���.�ŻFƔ���V	޼��2�p�R��qQ��;�#r,Z�X{��R�4,X��S��`�~�z`��)ON�J����0T��j�ϕ����+}���^���k����뱹�cs�?�1��]o��v�z��㈑�ͤ8��S��	s��_��
���T#8��M~��.wf�$�y��h�T�^�&a���U>_��i�o�%��]�߹�xzO���J�cf���%Jo{��"^�4Is��4y���嫂�D�U� �{#������A��ѨG���h�^ݞ �bJ�����a��x�XRk#��&��~�M���B�uʚ���/@��l�(|�{���#�d�KȵmD���AR6���wڌ*,@Eg:���V�����Ѭv�mqV)j�b��H�8���ˉ��^�ćL����"�1�$N� i�|�}/@�hܰ<�>��V�pH�ئU�̋� ���`�i"������58��b�zv)t�m9�'��G�����4ʳ^2f���0WR$t�wAT����4,�"��O޸xK"��>lS���X;�CQd�#n[y-�#�@�>V�cd�(�Π#�=�����>����;$�=/ ��PP��$�\��;�$�b�ru�Y�I��/�<��I'�1B�x�&��oɔǄ��N����	���_�����g(��@;"K,���X,K�N
�I������R��c+j����=f"��3u?��b�n�ٛ�����ڇ�*�`�w�5�~5@-,,��ir�K�mʹ+.�4�Z��1�FMR��U�U�}�
>�$a�ߤ�c}���R�A�~������ �75�̶e��܍��4�.�nכ�c�3e����"!�E\y\	UզC�%�Q�s����n5g���y!�m�Y�i�I�E%Ē9p%�w�Y��{�BjT�����}���?K�xm� v0:E�<�x�5kN���#6z��>��0)^L)u=�Q�m�k��E�l*�υc�Y~��f�J?�5^�uD��qt�-�i�}�S�=���;�����僘�����-�g���x ˔�W�;���g��b�P�mj�l�ˁ3l�"�����0ݞ����|����N�OޚE��V��5����W�V��¾�2KL�6��v���e���1!���Zu�E���x/O-CNi�� �A��S"���DR�͇d�;�
��d�8~�\G|�"V�B�6K�M \�Y;L���@(F��!�_��jӾ~�G��w7���@���e<� �.X��������]�m�5�W?n��h?�� �uW�v�%m_��6�,��M
�� F5��f��"��⑵���d�$& �Hr����iKU�������.|5T��5�N@;�G�d�����`��H�Kv�#���X�Z���9,V�2䣜���V�r��{mu�S��L<�5��v�RaJ����,�5z��,���9�P>�K�X�d#�m�kA�D�T4SQتp^�
Q�=���H�L�E4Z܉b��k:��˕�k�����u�2'�̘�G��K���*�䟎���}��:�<�y~:����Ҕ(�$�H�i�Dv��+[΋����o7��<Y���J��~�ċ����Dm1���������þ3�&��w�����Ԇu��m�Z��Ԭ�Dn�S'��u;@7�$i�d�?�MC��*���I hq`J�xz!�-hoF��L��"%2�P�������v8k�J�
��V�b�����´�X��s����^'K&`�O��ӃW�*�`b�j���W�d��6�߲�X �U�F��~G�@��ւ�؅�5,b���Z2�"؂�����i}}aN�f���\�s';����b���M��E/��GF�jE�+[_�S�Ͽ��g�i8��� $�F6/5�B<.�,r'M	~��V�10nG�]b��9�#�𲟼��l��V�(g�s�%XlxV64EB    fa00    2a30�Q*a���K7��GG��\{��+J҄l�Q��4�)/��wb؞��|���w�a�����bO\���(λ�?p^����eI T&6��+��'�FS�W�K���S'<d1�l�P)�=8\h��*i�3��.=�O��\?���n*�+~���e�M�X9$��i�Uü�k�M����dB��&�t#���1�P.Abq��&Z��ZV$Sw,�����	�?�1H��[�hy3����}��0ZI��7�-�=l�T�׏�;�{���j+o�%Uu��!�ޘ������bÑ�c	�~%k��9p�8���/?
�50��+��W	�[�ۙу�ˆ�L-�zu� ���]�:Q�TWu$��W��y�N�NY����U[�n��M�&v�MQ��;'��6k�`���
l=���j;˖p�V�ȝ���b�!Eկ*�0_m9�n-Ⳅ���H��$ ��'
}q����>�J���I��o�G�<0|C�K��[�ז�lSt?L�`�E$W0`����Ӈn��Bk�덉�����z�)<�8�$�m((�1;���4���������m��!�gŧ�2u� .׽�0Q)�P99#&��<��j��BI�J�sf��2��u#���d��f5�z�����uVr, �3���7��M�}�����\z(9�,v�'�絁W[y��s�ˋ@`�y�c���6�_�1��ʯrj)�E�b���ր�p*�t��	a<ym�q���O5*g�1��!#�
�Z�yOV"�/(UdV���t{��J0�s��A�/��ĳ�y[$:V ��}
.=1'���
�,hl��P3٨&�x�p�4*w���W�{�#c
8�>�<@�4m��+av���Dȍ&�_~����	Ʈ���C{3���N��	�g�G�+�Ą1�#r^f�L�����M-&��#œEu���m�bp@f�4矁U��-J� �i��� ��ps�	P��`�x���o_N�j;q�1�k)Ƙ�.�3�z�#��@F�
��3�~&�sN��2�&duj����o8;x��w�_f�;ܥ�N F6H��P9�G���Q�/]FXd2��:�~�kɼl;�GuJ�p��D�}�l�Ude�u�_
,
�#p�3�܃d#����r9�bde�cM�ߓ7�-i�=,!;��2{&Ly�R�h���R��vCqY j���bə�߈<��j���L1�פ:��2�4	a��#���HP�O\y����"v�w �=�'��g��-Y�����)�J�Cٙ2�mD��x�w�AK�n�������0*F�t�/��d�@�������P���` ����m�dދ����Na;l����K;�-�d�ƃ��@� ��VJ�|��x)�|�Iok�UbP��ivE�xy�&�i�����aLj[�7HS��¬��¬��Y�5l����7z}��X�.+��3��x��s��3�B��1$�f,??�~;���kk���{��t�������D����N��e�l"�Ċ$ C[&Gb��e���lE�Cv��	��
r�%��P9|-��s2Gx��3ܫGf!o���79��L��� ���ܞ�ؐ���hu�8}�
��Ub� "Eε����IT��0,PE��������k�� ��sfA�Z#>�?E^�n\H�yP��<  ���!��:�)>��%)o����&���Z 0��柾G&&W�Fu�&��`����hN=,�Sj���VH'��b<?��[��HV�L�5E�0��||,��)�q�kz_���ׇ'?b�Y��cġ�=9�M�[����,O�6ߎT��W�J�̈�qp���@T��(��EJ�B�T�PYM�|� <p+��+��E���1=�>b�҉�@���0"0@�M����RF��/��F�bB�Q�렶�su������>���a���ޝ}� ��4�!ըT��X�>\���e����I�{�0x$9�w�@�W�2ي&L�I�
�5�=Ǉp�[>���� %^�bV�s��V����s�,WL`�GL�UVo��<�UBO�J�#܌m<��v��o�7<^���6�S��Q����Ms����6�ɕ�{�~�Bv�#)�Dc�I)Pn�y|/Ј>j(ɖ���*e��i5k�I���[�v��<_�v�Vb�,L�}W|A����B,���6k�eW�{�����+W��n�K�Lu�*���%�n떾���mf���9�7|Wy�N�I��35�8 t`�$'�k���N%U���]�* ��Z$�����ܶs��l�LNJE!�yO
>=��Hp�U�!��+!cP�
�����!�C������� �rlq7	i�����|��֕�)�П�4f�$���/F��;�}yzHԌ~�T�T\(��/:�,���D�wľApP_�u�k����[}������o��5--I�.:���H'9��tp��5Gp}krm�Q�^��0�#�����(���胣Go�j$A�#�ȁ�Ls215)�I��+�:M�Ƀkѹ�^AJ��X�����h\�8E 9���Œ\�Ij(9�O����8n��lF"��P忬ę G�ş��hOC&5���`����C��'
�sg��BKjd=d`�KhѺ��{)�m	�3���G�j�N�S��νC(�:<��~�@�I�E���8���ou�&�yW��>��'����;���w�:�C����-N�YJ����F���2u�s�1�J4HA�n�����Vi.2���|��6d�)O�	|#I_�Ss��u;�-�X��<�DFsy}��� �_��x��	8�]���~�OR�δqM���CgW����#0q��0Kf�����������钓���"����y���F0gBoa�S��%ž_���0��s`G�\�2ڌ���)���͞D�C�섂�9���O��O�L�W�/P�X��9?��7;t�L|,�l�8¥C;�������R�}`p��GM!�NI�A�^s��V�P󞶂�T�Kf��ю���˷��+�'b@KJ�H�����F��S�ʽ�~]��Bs?@	/�R��0��#S[������}�U-�3����7I��u�]�Ty�����g��$����D��{���`G�JP?)Ǚqla���#�Yj\�7#
+��tߨ�2$U-h��1�D �����j�����`CP}痸�w]��)��-)����I���;��m�>�g/FU,.9�0}�iO�g�<3�I�� ��a�YQ�p%��h2���C�A�Du�[�cJ ?�n ��I�<b3������� S7|�)d�R��Elg?�G�_AwgZL�![D�7�$��4�U=��9�����(G����k��"8�>��o�,*��(
�g;
c��d0��V�'�aa��a�ǄI�֛��y�����n��nW�|�nǯq��KIq���l���O���n�g2���~E�f0�9q�����\C����Usz�/����u�:�1�B&��'$*�ق�Í9[��r@Q��	���X�-ai�e���ӴK,Ҝ��mj��fJ��=CH԰���CZ40���&�*�! ���9*^�{�aH� M4�w����~)?B�}_���6˩!fۏ��cNz!�jb_�)��!�V�ڟ�n�`2�P���v������f�XӞ����Z��8}UM��Ø��vi`Tg�O�U��W�C��xH2�F`���ĸت5��W͕��Iۂ��0*��>��J�_�/�?2U��9������S)�>r�ڈ�f�W!\���S�o�"R~׽"�K���^ ];d�lIN��6`?�r>l�F���mmsq�Ȋ�ʝZ�8N���`I�i��������;�L/h���̩�2��Z�Iv���H�g@>l�f�h�ı2�P�:v���U�gX[���5@�O!Їŀ
:�Y���$�᫅8����(F�ƾ�P`Z6m�� s ���Xz��"Fޱ�)�``�gP6Z&~�Qu!��֙��'<�+
���H���8n-��?��%p��o
9�uЋ�|����K�r8>>pe%|�N�a�l��G�s�j�3n\cI�������3�i����g�ʮVr`;�C�R"��@a��.�$4��W[��8�im'0�jU���N)Ȕ��.�?�n�� ��T����Rͳ���1��`��z����D(�f����c��,���x)M�u�%ɛ�?-�A�Y17�;Ks�_
ȁ�+�8����O7Y%c�n�kL*�ɜ�0�2�+,N�b�M;t�G@��t{�U��.�����c��Ɏ�CfN�h6Ea���P-��G*߁fh�(P��%��aU���C�&1Iq��|���'ph����q�m�x�m�G�I�|ο��ۙ�Dc5��n��Ҩ���Ye��y4Us����DHA݂@����3��^�
�qƽ���?�3N^A$%��A������_���8gM:�1PŽ|z �Rc������,�{�R�voX�b`ۜyc~�䌲y	i��3�/C�A�J#=h4�n��������QC����Vt] �\Z��w|;�ä�0�t�A���
)�!�넴�s���`�TD�ח�暥�n8�kV�o��sө�%K
YV�L�Y=�&̾X�����d��Ce��=�ˆB��6,���ܷ��s��Sa�O�HΛ������������:s���Ec�k�3=x8t��5�Ь��ځV��3��B���M�;u��Ͽ��Bd���]ڋ	TEUM��wz�Ri5iD�+��\�Nlk�"1>Nfo�577��y��}}�;�V��S8Z��H�CZp��>�v�$�y捬�gH6�-L�J*��b�����lI�54��M"���)5��	��-���q�*j\r��p�r1\`u��*0?,����\_s�>�o�)��.>.����[��h�;J˥�(��+�6��Q5�oj��2K���#��\(�v��?F�k5�@�؆����'r)��H���ކF�67}��T�y��˟zC�J��Fy+-b��w�l\��q}O�ʻ���^qB������$y[��SN��IJ|�������L��8m����o���ϻ]Z�=N#��z���w����I"ÈH��,��o�ɴ�l�5���G	��ObF�&Z�Ge�wȐ/�V��ȵj��E����	�����>��+�V�����#Iz��8`+2DyzF;i�?�˷{Z���&���]�G.)���ܩ�� �(߃4\��qr��;@�#�)[�Њ���J�kIߢ�]w��<,"�a�5�qu�����؈�EM��Pj�/b�:~���K
�}���-D������e{[��	-װ���}wdƫ�gnf[�x.�+��N:̵^oKn��=���ō�8�?�yӿ�Y^Қ����O��{����H���x�z��Em��C%g�5MV��QX<+�&�N[��?��o��)GU��]%?�̟��(NH�,�|�4k��|^Fގ[|&�]�"6O'�o[�K'��Z�_���R$��:�$,)�n,��~m_c��@�M'IU�-岌Z�J9���9�K�\�������T,�,���T#�̄Uc<���h��V��Ś�6��9[3CvRcC��X����Q�N��,ab�
2���kz�H�k!90�>��e0�uP��ה�����'o˷�9����������I�:��a/�>P��h:�=�Gh�/�>א���Vx�HR-q�he�2���ûo�9<ko����a��I8w�&�R�I���^�ƌB-�U.IA�� 2[t)_���%�
�$�V~��oo��b��<45��8-�����-�YZ�dt���6��G��Em�GD�5]C�r����US?N�h� �8L��]c*q�u]�+ݢ!��� v\�/����6S�A��H[�_� ��4F=���v�{�3P��G�a�pu���,Wm���dBA%e�E��T�{:���ܪ
�P5�I�ze�x�a|�g�
չCN;���.��z�?�ڬ�Ma\8p&>�H��sl�Ν��L�H�@v���&Ӆh�U�Q�It�kr�o�4�l�>��Kָ��o����S���{�\��4��˼�rd3���Jc6Y )D��ڡ�@�ɽ��e C�ep"�!=`��H�-���e�iG���ٞ������N
lO��s�HĊ�Q����H�:�\�-Ә6��.�)C�q1H�	rpz�\͑AH���lgP�io�Q�~5�d�xvd�&W<s܏�����b�k?�
Y�n��|��4�ز$
|��,ܰ���_��/0���	�}�Tj/������)�J9称 }K���})��{I���|���)&lJ����)�Wѱ�"۔A5��6����k0�*�WH�T&r��2�&u�C�[���%�YeSp\� ��6IS�ැ;�W7���@'[�	R��{�e8cC��v���ј����RWNȊER;|��V�~����P`�[�l�t�n���>�s:������לn�1����X�ٷ|+�r�G�P��y��,j�]�?�Q}�>�J��f��-��Z��/�f��Z�^��(_�[�Ҧ�ԕ�[�Rg�< �;�#����DM쿌a�Jik��6�}�eQ����o�[�g�.'���ŵ�j/�D�C�V��%���*��I�����u�-�B-/?6�(�Dm����k�^K�F�д�����<�5n&C�CCe�On�sٖDz��u�?��Hj�A �=��i&��n"�5,w�,�8�5\���'G*F�)>]#��7�����3�Z�8�@������}��_��N\���p���)�(�[H���+�X��~��d�V�ߘ&�!��x�8U�r�� ު4̨�Dߺ���N��XnVP�Z��L��Kc:�-���*��<���L1��h�H��t%@`�g cN��Խ�k^}�>���l�8������SiM����44�}���#;W-y��J������)���w��l�o$��*n�ECeĳ�ؤ�?�醗Z��:���F�ņ0p���B�Z�ϯE��7�q���+�Jy|u!O��G�=�8�Ch� W�M��	���1�
��!D�f$�᪌w�n�B�^(Q�8E�"X^z/��R�� �����%���<�D���x?c}�5�"!^N��wx����QtV�Bn��L���c*cK��g~]���C��X�=4v���n��$�����*YY,�wg�&�峇��D��O
�2�;�p�.��56�@%b�)�߼�+��Ӽ�.�:�<�-v��8�1I`���i"'�OC����Z|��_�~䴴���OU
��Z�i���slP�$�VGM�V��zi�h���Dc|	;IuN�g���-7��y�x�:&-9��2P=��l*5�G��&�kډ<��Y?��c	�SPmKJO[�HZH�~>kF���Vi�Ή&�ъ*�&�����*D1�Jߨ�rd`�@\�����z���8Лϓ��k�!���f~�Ka�=�n�f�K���5�9?�&��dq�!�-��Θ�u�ГC2�OewR���a�u2��B�+=���t`��*n���Rѫ������8q�j_�aVn�����}2�$ ��B���4P7��3߭�ϻtf �G�([�	�	7�bn����C}��E�8��
�����c�-�7��x3��R�r������Y��ڶR.�j$G�����S-,�CE(4(m��  /*4����4K�mF��M"�-�F������9�
ȟ@e*؏�7��|���w�B����j4�Y�k�<G,F�
�rΈW��yB�����n�[Z�ܴ�ϓ����U�ku*F��!���A�)�k�vo=]�-�A�Ƅ� U�2����*�%���q/*]M��~3�!Jh����r����m� ���d������i�l�n������\�����A�׸y��ʗ*�$>/�H�!�[��+ݲ�6�]h��5�b��L	�9#�����L�Pw�#����Hy�8������.�<�:��oo�_[����l32d�p��:� �?��d�B*�{�:edt� ��&��09	��^�����A}qmt/(lH&�*3�Z�R�]I6a�L�j���1'���o��X9`0S,��n��oF�ߥ}�A��a\ɦ�D48m4aYC����+�U��z�/��\)i��_"���o�D.�Sx�b��oB�	wQ \t�cU��g���~�m��3":��T4 ف19���r3�����<E�]��Ht)�>��jJ}�b��}�M�2��? ��W@�U����^vy#�)ͱ��Y�^�鍧rǩ����.�6-�5�Y�!O~�C����j�R	��"��3���\�,h7b�����b9݆���i~/|����]���,i��y��3�N�j�K�.�y�N1��f@�ݭ|��cyfVn��j�	���^b��Uf!'���������m����gf�8�M�E���$��+�c���K��=M�Y�Ԙ O	60)��D^_�ѵu��KTy�((H��j&��M���8/h��Rg���\���H � �1C��P���
����}�v��R��c2�϶�T"{�
"���F
����Qx'1�]���^�C�<��T�e�R�6ǀ��pp-�q5� ���?Z�T��=����B��H�*���#��������Mu��&���'��R��7�g�E>}�E�t�j�� ���Ѩ��z�?�G1�^��U�?��
s+�V�i����2@��Qa��P����k�����9�2�R>�_���5��J���0�"=u�Ջ|Z��/�f�F-�{Ex�od[������C�N�-<k?��э�m�)����C�\�$Ң�W6��?�����]T��v>n���%� ��f��uC��0�=e�&G��B�8X��a��G7_��b��#r�x/��cG�5���9����έ	�cWs�pd�lA:��i"�yr;�&\Fn��v�5q��q[Eʈ�?�,p��ǚ�Xm�������������A%�B��}���9��#- ��=%�#*0����Z���~t�	���j B4B:���-㸱�l��P�ZHP��E�O��__�A�h�|ǭ��\�`���D_[�,��tL0(;���������4�t�yr����Յ��Ra9����N��e.�����#�(�K�0�-m��N�Up/�LD���������P��!Ҫ���{�LF�.y<�a?L�!�MpG�:,˻� :�!yT��f�J��C����P�q8-}��<���h0x��;X3�k�TsHˠqLunw�a[(I�.��������*�ּ��f��H|(R��]B��q��!̔���g��r�{�GHI��W~�h��� ��b�T��f)�;V�գ�)���+Ҥ��	5������)�������m��.����`a��cGx��Rv�%�V̙������b2�`Ic��Ҭ�*PJ����s2a5O�>�
��Y,/��3y���UK�ٍ9���-������#m����$��n���1��αI���Mr�@ǵS�q��"�|��i/n��Ui�� ׃���pQ���@��w٬��Ev���
֚�y= r�<?}�F�/RP����2��H�hVM��|�F��7���R���3:�����P崝��h�M��wE�sERm#�wU�dE���zLC�{�X��S�g���bf���[1�rL��ژfu������c�M9��w��W^�熯��Ę�AR/�9��U�1���ى��t�ģ�wam�<?H<���J������.CV���]�'\|�&T,����w��x��9��E~gb/p�,y$��K?U���_�h�c�'�Y��
B��i�ߘ��
���[��A$jXGy�����P��W��
˽����i�K����&�=�{��Iw�qm�E,��W�_�j���J��1�zS:W�r1۪�2���RXݲ����������ޒ�����7�r'v��r�V�ʣ�&��|y`�V0)�[��� �uz�.�ՠgt�yK��f�� �>o�4
P�p��[��0(�T)(�T�0Z�!���G�I�P�=U�@֯�\�k�綃����+&s�U�0`��q/����g�g?�
]�Pj�4|��gU�1`H��+E�"i��S?���l�"����؍"�9.�
R/�z}��ʾ��pǈB�43��gB$%�1��6]��������bb�Y��.� �KM�b����<=�-a�c�+|P��g������v����7�������X�SQ�d�^�J���%1y�s�	&Bui�]ő�ŌD����mS��;��s��:@s3�������z�҃�Rx� "������؅�Zj��f<��c�qa ��q"b$��=����]�W����Q�Y0$�h��'Gs��0cӕ8��'��5x%��8�"�ߝ�}k��5���̨�bN�T�O�e�Bs�.5����l�w;�a��&�ϻ#���]J�`�ef���VL�YU�b��nM�G�@\z�(N@��u�M��&`#it9��Znm�s����{�����'��T��ի }�D��h��/]}2s5���"`XlxV64EB    6053    1320T}}$VB~�jE�v8h*t5��i�QYb"4oǓ=O�U95э����Cjb�[Ў��'�n.J���va2�	���+vc��r*-뗄r�!���}�A�-�t�Ab����0"Eo�XR�D�I�K��ڀ�����R� lE�Vg ����(�w����K;���I�:��PJ�ŪW�+*�id.�K�ͫ��'�]Hɷ@�?�5������Xc� ��+���3Az/
���w��T��T�WPh�R�5��'������Ð�6�a.{�5�V�|6P����L���L]&���>��������-B���ih���0H�������eO��'7n����ݍ}o�oL��j�g-t�ʝ.�F���Jfu<��R;�����U�ٍ"�cB��bq�a� �Y�3�G�E��P�+������	�)�2�w�g<������� ��YG��sH�,��<]�lH�G!>@iq��
:���2�o'�֫
FjA�o�.)#���ׅr��΀g���V�ݠ�3��Ďtz9P��?��m��F~�i|��ݶXWC�
-ǀ��wZ �T�b���M=�5�6����h�'��-f�x"��`��D:��؆-Y�7��A^��踙�u����۟u�R[Zt�b���W��sߋ���w|�<e���ux."��R!o�k�8�U��f
����/?����k�G��8��K�Y,~\��w�JPV��������U�R�rD t<w(۬/k�歅A�0�"����SP�k��hB�V���#�~�r8~����[���K�՞ �RU�ũ�o�4c��@�a�w���ٞ�����J����&Q�Nr.�#w���7�-�=>_g��V����F[����8Ti��պ~���vܝ�<0-�ڼL;<��=���u�s��g�Co�1�U����z�ʌ��p=��W�?�8����F�w���*m'R*Pb���^z>] �#|�Ĳ�r]��#��4�G�@��"31�8QzN�3p��b��-OZt� ����;��"k���&{�UV��Μ�MH9b !�*fD��Z ���2�6L>v����A�S����㘂Xw�A]듮�Ҹ�K��\�g�S6~���!���va8��WiK�-~k��b�B�8���ƌD��W��φ�	�B���8�9<�I^����0k��0gk��Zp �ir��� zyt�u���%����j��	g�H��&J�z4��֌k���Ș���ɕ������+eւK��JmD�^�PSl9�����Q2a�\"��=F7$��.��X^dWe�c��d��I��W���C��~"W{�O+@j%��̳�ܰT�X�]��>�}����ah���_o����q$X-rf� �v3.?/K-}a����ߥfN����(�`��i�j����qg���E�V8#z]��r9��:H�>�i)�8d���*]�7�(j�)? �^R��Acƕ�/�^X�˴=�S~_��� ]�b|	�=0�y��"vb*5�6�r��J�ӟ�O2�%:>�`^�U˂�ל`��}�_�B�·���8O����04lo> ���STO�H��Iܳǻw)��*�8�i��2�%����
>��E�Ơ��T��[`7	�����2����J���i`,Y?V����]����{��I���x����!T<�ϸ_V�^��I�,iy�mU�zI����I�&y��k_a=ҿ���s^f�[Bq}�驓�@��>���B��)�)���cn"�*�N;i �����J��*&\�ͦ��<�wvF�
Hz�����wi�Հ��QV��VI�����IFg���W�ayLZ�N��%T@$�;jS��V��'�*wBG����I+qc���څ%
0��R��.Q��$���5��QQ���G�Я1��7k���5�N������?�'��̦�����/�T�AҡÆ��ƾ��gk/C�l�?Uu�WP��ݔ5ؔ��x��Ѷ�W�+A�� ��
���։�<j�V���q#Χ���G�wB� ���-�=W�r\'��\Xi���?P�D���n�73oQo���Y��~�3�,#��MD�/���M֖on3�)�*)�g�H�z�ٗ΅K�cvؗ[����t�4wϩ�W���aފ�۩ڔŊ���~�V�|P ���t=�p�#�
8=�������#G�Gr���è$�CrE�� #`VN|ȋNˆi��P�1�N8>�Q���=�3?]薃t��U��Ȟ!�>�XL����o�
D��%�3)��:һ�=%�Ho0h��*��+�4N��0|��y��xx��Q10BǷ;As0-������_%=4�-A?�MڜkDYh�J�s1�1��r�
ɽBX�7X23o�N��������_����v�Y�%�ڮ��eoT�PϷ��|�(ER1�E���`�m�s����Q�_B����D���G�|����V���X���P�+oA2+�F
�)�N8�t��=�ψ�P�Ly���2� �]��%6|ԉ9	[W�=h$��9�m��q-�%*�s
��k��e\�����5��6��T��d8�����_h Kz�8�)gw�sf�y�fW

(b�]«Z��9W��y"3��0w�8��� ���2�D��CC��,�.�<���h��e�d�r }#M����Q��2�(tt��dB_(/�O��Ǜ�s�W���Q�n�2�0�� t<�4�!.`��s�{���on�@J4��	��Y)��t\�ZRf�
E� >��4�a���S��.Fp��1vz=����IDu�㓅,��.�5d��,Ճ�%b��U��~�6/��3��G\�[eoL��Yp[��j�(UB.�mq�'/^�r~�*���n�+'�.��v��u`��A�F�~[���w�3,{у�Yb'<�;2e�:E�w�-�f�.�$����A%6�^C�I7%K�g�ҟ5/�!.1A�T��6>��\�
}�>&eh���W"�G`���e��-�S٠񷷏#�:���=:��槣��h{����x/+�W"���y&�S3����!�)W�b�p�XL�� ��aږ��?�����W~�*�1_��t�$�������tUH�|O�� QD2��M�ݘ����ڌ��/�����^�w�^ṇ�o9,G;�朹��a�����\�)A�&[�O�J��M�{<Q�n����K���k��o��I/�@��	�����,�0Ա��:�%�'4K>�(�$k9>����6��aiy�i-�O�to�����i�P�L�c�%�z3 �,�;Kt������_u�R![3o�󜢒��XO<�����r<�W�dG FK%`��=8���������Ԟ�k;6��|o���sh�D���|XL̺+p~�~^q�	�6��pWd�_�B�8C��� Ɗ�k��r���� a�sT�!�7 ���#&�(�N�m��S �㓆�=^�MA�J�t�������iƑ�#���6�@���@{�mE3�x_R[�[0�ߺo�P�w�3jC��[�=F�f�����Jf�9�Y��a��7�)�T�C��&�ʆ&�hܔE��rt�r�"I���{��<��f1�Ϧ�L���ïĉ
&��)�[d��K�?�y�/uÀm�A'��f������F��t�K_�AJ�KW����ہo���$�Ǖi�v���vQ�`�h�řU;t 	Qqq�t�?|rYH �eK�Z��oUUDn��#�n� <
}	�(�G9����|u�T���j�w3�O�����u�����V�t͛�ޅ�����d$�T|"���.�rʄAh��������MՆ�c.����_��H�����Y�{	pC��~cQ���� ������� 7b�؊c*l��k���}�W�ܾ�,G����u�;�A~-�
\(�+���/yÄ>������?���jl,q�Ł��U���ϫ�l�9����{헊�ش�)K�4��"[��j�
�D�8a]9̛V�Y�O�yUB���-jf���mt��l��٩0��@/5;�th>Vt��qe�|G7�0����&x*7^�~�)k;=�&���BG�}pBڑ�kNÆ^�л��9o��6��#R�rMnq��X��\BԨ1x�C}�WC���^\64���4���Xk�Al�͗��ױ�����!XW��*da�"�Q�w�DI�rPX�������p��������0�:'���)���J�߿���&b�.s>�x���^��j>q�:�dټ-[퍜"3�7��Z�F~�ٚ�8�@��o���Zkh��˺$�B�����;S��0��_��F=ʄ(�k�p�\��s����c��m��$��B�(�C���j�
R��f�'�|�V`�4~,����
^�m�/÷!���#L 2���Aj��<W6�^Z�,~�BDAh؃I����&�-��d�H���^�V�Db�g�Ƌ�����ڃV�lwg��A8��,)FO'����~�������2��[PS�^�(90	ney�AE#��z��'�`XI�� T��U��`�Fmkc	��_�/�`K�vF������!��2�12t��A��f��L������jո��n���@h�<3ȉ9�8�$�R|<{j�<T,�#�ן���l�'�~!y�]�P���B�骟���K⯠�$xr��K])�[��v7w
8�ތS4b���/Yg]���ʦ�;*�;Y5w�X�@#����R���
��j�}�7oU�]#ڈ���ʦ�mV��s�xI��2Z�