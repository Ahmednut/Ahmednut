XlxV64EB    fa00    2c20�-
��$R��	�ј-ǥ0O%��n{s�����΅G�>ʟk��*&D࿚����{�PL��c)xt�
�""�Ȇ}mm�`�~>��˅����ؠxL�j�=q��N��p?�0qA��TW콵`1���"g��<}�c%��,��g���n,}�	���o7M�~mH��hY��n�7���6�♇��H}ն��pY2~�C�lḚQؾ�����xg��iw[�X�_}�اH����-\�~�ט�e��l&Hy��[�j���"�����6��ޣQ� �u�O��aVq��p�(�P
����j�-_1K�Ps׀�G�B�~���j��5/��{Сý&>����zV;6Ö.m������-�����y�B�sra��kW����:�OOQPxl��6�WWRO9�h��κ���w�Y�]
M]�wH� ��PޑGB߃R�v�=Y�+�� -خ���D�J�v3�t|%������ޏ^������'�4�՗�D������}m 
��2���tԞue��V ͢y�UM�5��=��M��Q��A�a��j����O�O�OI>�I�o���:�*��{��]��.��T��w���Z}�����d͢\�Yiw"�}�qX��k�[��|�[�p�� E4e�\���x����B-�$����d����~<�r'N����yg�fZ.�����q5�r8�`��E�T�2���P�vIK��'�9l7v��G	���E��?�O寑�%����ҎU�H8�lh�����d�	�%�(���_�׸�֑a�w�ʦ�\+4�:�[�8�����>�>ZByO�'�햷�fy�{�J��4+�2�ڙV�	}u����5�PMTE0~��]�Qz�(��ġ����h?ݷ�^�+(�t��_)%����M���qv��״b������#R]��f��*���EOn��5Q�e��!����Y�QS�߶���f�k�{
 �j����4�Jl�L�N�����
1A�a�������Pb�,�51j2J��rv�*t�j��%��˶q�����]δ7	��*ϛ���d�/��|(�j�$��M�M�.
d�G�Fl��.����n)�@#���9���3���ٖ#hෛvzl���-J��H���'�\˝�7��-�,ǟ�V�l�eeg�ޔD5��s2�2�_��d%ǃ������][��#�(`C$��^O�H�E�(����6�gQ!�߬�`f
sə��2Q�F^�Ơ�k��\%���
~�ܲ�u�����9E�M���j�lx��%���7�&�ج"����J	�$B �����$�O�����ʺ/B��2�n<��Vk�0R��Ǭ�oj�]�U'N݇�d�(���v_̲��wpŋ󑿶z�H	��2�	���@�M�00�5ni���Vs;<��x����@T~���g@��8SA(�&h�0@�b>�`*)���^8��������^b������:�g�Wx*�c�	 ����9�%������-�/M�q��q�%�d����_��ڹ�yS�&q���J-�2���K`�Q(:g�d�K�YV�]P �4��A	�]�JC:�K՗�mط���̟�]Ok��k �Iê��~y������	�-+A$5��KԿ7М�K��4�PJ:l��l�`f�޶W���~Kz\)0C��W$�/k+��HN����q�ȃ� %*�Q7�8H,O�2���_����̻lφ4���a5�3���/�.v_
>�ē��;��%&�`R͏ED��\+��:&R��YCK��a�ed�}��?)�?��ԃ_IӅP�yi>��$O$�࠿	ם?(��g.O�W:�	��a3���	�m3"2Uds�����G�o)���7�dD~�����h��j�$�l�˜
/4�!�i�0AXK߼����~k��ԦM���{�r:�n�ȿ#\�85w���!����6N�� ۛo7̊�%ZBF8�5�my{�"0*	��3DwBy�I7u��k�$H&^h�bk؛��!/5� -��@)�����e���R��|tS4�ఽf��$��2����[w�~u�Z�$�ڦ}�O�A��Hl<�Y�c������O���d	[�p��<{T�F3�
4�ϑ�/s3$�*��H�[0���c0��U�d'�	�KFm�U�M�?q��r��W����ެ>�E�J��hp�]~��Yטw\�������!�͝ ����I��D�Zawp@z$�Q�n�.kO���c�
l���nC�=��~�u� �/��{���S{%?�l*��B�;��ZX}R4BB�sz(`#G�)�b|8l��Y���������a(~Ε�õ�峢���������}*��J��	G�g��eZ��3j�m��UJ��j�(�+��qDt�t�m�[�A��|ɋd�yP��0G�6��o�m��h�դ]a�O��f�7#���S�dhĝ���5�?|Y"5(]ʀ���$tW_`U ��{�v8Za�&b�M�Y~�P�n�0�3w��M�Md���8���h�4y�E��۶���`�I���F�
��R;x������	7��{X0�<�����|y��18W�m��S�~�Y�N�他�"��e��Cw[$Y����u��֧; mh0\w	�ֺ
���e Fx���2����)X�a�k�u�\��D���~�g�B��>�@����MC��9���M6�ͥۧGh�yg�3uwF᭔��Y�57���e��I��i�t]<)Y5�`��2�E s3��1�u�m���8*R��M���f7f�%��!0�e�j��U]lLJ\'�h0�)@��?:1�tD m��ڎ��1JL$�akt�?��j�Y��JfY�����"��q�#p��7� ��G��M8�g�����$nb�vv��#�=�����d�;�炤��!A��Cr��9�8���� ��Z�������$��� MP���
"��V-DX�����O$�H��ꅥ�|��^Lu�뮬k(�/m��a?O>�6�I���7BI��[��ܺ>�	���Tf94/J)�����S�rz�z�>�|�MCJ�HU����@<�wՀL�����+����#+D���:�r@���	@Wb���:�gM��z��4�
ٌ���V)9s�:N����i�ד������9o ��4����I�y��K �yx��r�x��b��+ѻn����
����ˌtH���C 
�.lw8���{�v�ǃn�<H3��&�ύִ�2��0�'	������3%�?屵��C��HO��6�1��1�}�+�a�^����Ě�K����,X Q��mb:d7�e���� 	чx4��n���k L�ؒ|l�B��^��7e|��L���y$���.,���rm����k��\K$U��@��S�x�PS�,��ʎ�p��f�Xq������Ȣ��'�
�n���l�����e�Jm:�e����t��@��
 �3�^)Oz"�ك��!�E�'oҁ~�o,��)�Iϔ��A�	f����C������4��?���t]�krN�r8O^ƚB$�c��[�^1Ѷ�j���p�&a����&��}�������5(k���{�>�� ��(� �d���{7��\��i� ������֋͐��C��~ �c�����$M��C4��"#���-^*Q�G��� �j�4��kĢR5*��K]}yY�����	�u�}V�v����Y�92_��o�L�üa���#U��cfj'�u�}$� �\o�`~l#�g>Bw@�w��dzF��$D�X(���K}"ap_�3˯�){ ��C��i�K�Fz9���jv�odbe�� Σ��t�!r'�X.�=g�~�k��/�����ἄ5WV��B�>��~N�2J���'K���������9��F�( E8<9��ִ�Pg�T�*�f�v��N0`�o賰��n��>w&5ge,E�9V�r�K�N?�%�M��(�v̷	Nm�]g|��hN��w#�U�H���tT�Wz���|�G�^8���XB��$�5�]æ�� `��������k3w�����!��	����%�x.&��Ҙ�x�Gi"��������$A����~~���5�֞��5�{Ў��e��*S���oM
b�63^)$��K�H�+1P㎊L�?#�A��s���5�j
`����y����r�����z'`�w��T��θ��"��A�
F��aIq|���	��K��$�p�g�ѣ���O��~�6YX��E\��D���V>�p%��
@,A��@#vA�
a���tD�p�3��c�{8����Ҧ?���9B�01oٙ�*�0�	y�䈮!�Ԩ�.��X#��K�����AgB��XG�"�h��#[��l�(e92"�ClLB<���[t������r2k���͆3DT��nG���y����+����3fG���v�� (,L�'��bز�jHRoi�x�B����
gQ�Cs�}v� ��E���0f�}c���M�޼B[�*�Ds�rO$��_W���W�?|�� fws�~��;�}�)�^�\�бc�!�\6@b�e���$�T���̀���i6�ݕ�ݕ!彣共�;�q���N1T���@��nH>��8Z�(/ւv6>=~0�On�x��f���g�=l�шP�7B �;�0/6�����zAO(�8���>�Ȉ%����:X{�<���V���y$�D쯃
�(\nw��K�J�[+�m�Ņ��6�����|��=%�m���$S�F����tL]�U��q;k*<;A����9�U��"����*�9�ꤨ�+sV:1X]�F�E(������s�	O����2�9�i��g3'���Y�:il�nh%}2���_��G%��;�H�E8:^��q�wEd�����5����ǒ�2���Qc���Tv�Xxx�c�$(�Y��z�_!� �9Ŗ�B2h�ew��<x�Ie�Ÿ��?�ۇ(��� �s�S���ͭ�!��J�!�H,X7�gC�]��`�w'o{s���E���0��h�^-�@ �:�Q��i/��s�Fm��!Ԃ���-ޘP귖o�V��L"��
���!큤H�bOn��1���Ax��0BR}�8�/���e?�(���{خ�a���mU�>�A�9��~��|����ܺ�>H��Y~����O�hQ8��y(c1�Ye/v5��|\`]��I�X#�e*��  E�4ҍ�C'M[�	�Ch������	�D�d9p�������{^�t�aKO��|��rCX;mBav�gv�&`*9��fN]c�V���⃙5��J�S
�i	�y4�j�#l��u�Sι�Mm�ʐ�'a���l(�0��b�
�3<=��A�S��d}."��~a�,�]�M�!rt�W����n�܍
k�Wl�Tc��H��`���
:�Lq`8�A^�-w#/�'��A&FAhZ�I����?��3�R��� �#W��w������):��
<q�j�|�������"M�
��m�`%�uD���WcWǍ%�2/��z�s��}��Ǿ�Ab!�������ʮQ��F٥��W��p���X��v���pna���e\4|OqլW1���#�+�R���.d>7t�D��!���MT��/����}kwq��g_B����Dv��{�(�,�bY�~9n ��]�TS-h���	���%�޲�F�ّ�3(
�'�O} o,v5�ZJD��H�ɒ��M�+��ΜxU���'֙$�<H�R�f[<��
K?&\�3�{�4o��|R{���MI�J"�NΏ\rV��>�nW6�	��2�#y�(���N�g�n��A�V7'���"|�F�����r�#1����f�bSb��ۑ��#�{5�Y�'��]oN��l@��4�Ttsu����iQ���������gi:œ2�Em��q�~T_��Z}H�l�>���=����|���$�����7g�
��5��d�i���m�sb����u?��mL������s���2��@��m[ͷ&0���]Z�$��F��ɹ)��?i�7�_�pB�g�����r����+��.4���j�iq��B�v\J���?C<�n�,MX>@2^�ԗ�bl	��Mн; @ tmd�c.Ѥ�[�ҷ��L�����V�(H�q���I@ݞ�t�_��k벺PX�X�|�P��$���<���y��[\������V�\o�n� P�d8z����<�Ο�m���Ỻ���\�ٜ�>�z��2מ��5�������F�XH0��Ol��r}�C���k墘��?�(�7ӊ�9;|Zk F:U5�����ҵ:�D�������I[ޛ�k��lW�}��)NMi3�H-΢�kc1����m��meD���W=	Vb~�j��?�1���-�a�7�5:Gr{w�t�:q�ū}���$�b��{#A��F0j
��#X�Q���=	�8V1�YB_���i��4x\a�cb�G�} �Z��V�⯖�4�0҄>zk�i�˖�g]0�k\�4'�8��@8@1�wz��߲�̧otk�9Ll|�: $��o������Yz�t9���r�P����K)�\�\�Kl�n���Z���@]����@�0�^]�K=Y�ݡ�Ԇ��g�R�v%i�]L][,�3�)�d:��ų�A>��%~�����A3�^&?��A�B�ɠ�83�\��	�qإ�I�R�eRe�I��G�g�i�]X�V�{���f� /G��װ3V>9Zu��n2ƽf9xkMվ�E���^�z�ҒNDJ�T;a�28�h��
"���~�$�;Y{���p����Ɔ��wW�9�3t"����%��k�${����u���M�����>3���`p|�`��<SE1���Q=�lr��ݾ��]?	w�J�e7E�h9u�<��m�e��p8RH��$�-=sk �g>��tN�6�1 I0�Jɀ�K�T��_^�-����!�����V�g� ��`�kN�!��{�m��˖�4lFE� ��N�k2��_*�����D�K�Z�qe� �ˁ^Hz�|?�k�x~�A���[�\ʛ�y"�ko�ф#*U�8�j��S}�_���/Ǡ�)���L8��N���;42���b�x�"�?~�WqP�Q!*�	)~��dZ
�Y�؎�eԆʇ��7��g�K	÷���UU��ŞK���ӱ�{?f'���ǀI�aײ>�;
�N`x�x�t�Y?������[7��-��0�ٞ�*[��2¿ބ�e-Q���V�X����`���1�P��NH#-Uժz�����`q!��Yˡ��Sv�X�T��[
h>��	���Q�����X�X�?��P�"
���;k�[��/�և���&i��dC��H��\XO5FDܸw����fqԃKw�j<U���'���5<�bD����&�
�ԭ@��J.�[5|T���5!o]D�_��}g��m�b���S���U����cZ�t�|��\�iRO���9	l%k�y�\�I�a�fx�M��,6a�D��fY�f�"�<��:
fA b�dU��1�7�^P�3�\�O�߼����z���צ����ɫ�
�� G�$���>���J*��̦[�Z������-�iײNx���[ͻ�/�?�֔X��o�P���z��+sz�_�0c�0#��\�k��n �T*(��B-w�3��MA���8/Q��}n�������X�1�f���2���h� p^�#����MV�n
�(mr�g�F%3�7�-wyN}�i"���e�FE�k�l��2Qe�wc�s�/^`�4-�T������z��,�.�i��B���C>ƌ������W�S�w¼K9)������`�;��U�a�-�-���dq��zC�yF���Y���>z��'�Y���k|�w�Aġޚ�wEi��;Ɠ���IŻ)�����>!��&O`ar��ܜE��"�$�+��'L�+d��b�$\,'yn�Bދ��+�bi��
�T���w������v�ɨg��t�t<670�uPFK��z�d�%zتʧ5
�H�$�ҏG�n��*�@�8"=��k' �y_���,��,�2�>����6�H�����i�i��Q�~��1R(db��:-ڌ��&��JO�)��zo��2��?c���We�0��>_� ����F��C$I���p�s�V͑G:�S LM%tِ��RF�[�ڬ���xǄ�@�=wRd�uX�n������4ʫ���*��e5[�ؒ%]�g6�T�@'�uyX�rK$�{ q>�iZ5,-�������;;���TG��}�
��:gJ͘RQ�8�hs�{ڰu�Z�4����µ=���o��D�E�N�*���ƒ�mɵ�; "�l���T��w���GHu�_E%Y���!�r�8��T՞�V(���}�B��;�V�&qa\�s�P(\`��"�v.4�8'��H�g����(���s��,}.]��T��E:��|q4�d�ų�{�=-�d����V��V捀�v5�f�Br!�\1�Ȃ�V�$^�^�W�b!�A�+�������NlCbߊ@����r'������ ���;\a��=��TKq؜mC�G�����˦�UyDLl���y+@��74��	*Ԡ�s{���F̳�2�i�NN/�*��t)�x&�y��E�K�a�y�8޾��g�b�;/`��R��J�h$(I'5��\D�%W�CBKJ�,՞"�����WWn4��B?�2GK(QQ�q�$$SrjWh�v��,���"	B
H�Y{̣�s�
q��G�iϺz�Ն^,k�Jڽ����3,>)�r&��=nfʯC�I�J��0��)C��y+�U����I��`�!�z���N���[h�,��<JP�y���X*�����k���!rC�7�5-(���_!��|y�X1i�ЮƼͣ.㍐�<p\uH0��V�_�u$+�:W_[�C���؝\�u�Z�:�c�v�X&j����@��~��\�y���ֻX�~Q?t����_���H����+E��7�W����g�����h�&V�C+�������`�k��J��N󲰡k�	P�g7���c�Uט�N2'�Ǌ�����V�!�f����@w=�	hY�aJ�!�*�yl�'I��Mb���S�ؕ�1��`Ir�_Db,��]d4*vI�;���U;x.���1�����'�8��U���smܴ�ls�!�ܚ��� !�\������pyI0R986`��
�2~b�UGJ�]�B���Y��{����)� ��&#uD#(s�Nf�V��[Y�{:��}�o��Nhv��&����~��mg�ʹ�YK�=��c��|1��� �sM�BA (m쓘�����&���0�J�U��8N���\ĳ�D6�����B�w&�b�����J�Qp�A�H>V;Q�����rnv�΀������$�D��)�J5��0Xx�?�9�B�l�Mh���0*��E�����
��������e��+pd`�Tl"���Sz�a}�2�����)��,d6tF�
;@Q��'�a�8�CK����G3��Y�uC6C&���-݆U��T�����?����*'��Τ~�t�,Y���bC��6�3�u4��t�.y�7�JQ�t;��h5ΰw��v+�C���-V��J��r{/��2"^���J����j�u _�-�K2�o�&�3qW�Ͳ96���G�l���p6��2�p��K�^ţR�И؜�d.�@w��vܗZ��K�ώB���P�}�IO2�2���k�HUL���Aˬ�ۼ(EyDZ���|%�Q9� �L�q:�'� (n�	���huLk+?v8�M7�3�21���ܣM����;dj&�JG� `�\{Q4���P�|��:��Z�Pz�y�W>��v��w��A��ح��p��dů�a�1AM��^�uod��u��m��33���i�IJ�;�=��1���2Q������oHB@0�����'�����2��K���Q7�]�b`��Pҵ�z-��D�&�.��6��:0#nި��&P��!{��t��d���e�U-�eA��̗K!�Vo�v��Q���W���R���S���p0/������&eN�5�휯��|X~N�tF�c\S� ��u���&	��IhS��S�y*S<� k���&�0��j�}?�Տ�^E������f��k��L�AJ.
&�L��槀���F*�7���"XU�(��2[܉?��=��S�@玤�l��ۻ��H��3�Xu����)]��$����m[�rb]:d�/��������%�77�B�`�#����=$�A����"�`�F]��\�?��$�\W��4�Rv:��i}ת���<L�� v�"5jC�|��)�dE���uO�<�I��(��LǪ�]wR���=� y���g��"j�K7�sw�NһI��'ؕ�O�XI�u����emP�2J�:�Ŝ.a`�@�Pю)�4��<�(�[�op�(|/Ƶw�rR� 3��i�4�..._�Vuye��nPB5�e���(��{kƸ7`"@@��Ɗ�|w�y `l�Л�Qe%�C3n�a���v���P#�fn3�ȯJ#L� L*�:lU3z��0�����й�6�u��R���f&p���DJ9l�W�bA,ɵ)MAK ��	����q�� \�rK��Z�E!o����Ï��*Ѻf�0 �Af��	�:v]�zO w��j�(�T:F�T4��i���R�[{�~��&7�ma�5�)u+���%kL�n�J��Ug�g�4	\��Y���U<�����|ĸ$-`�H��9s�诞ptӏtJ��J��ܱjz\%�|�R��@����w��(7�b�o6�����u�|��Իzy>���"TG���"�b���-+���) ʾ�~��ߛ�'�j�<�]�k���#r�UGmP���Q�7��1�{	TM{��4?A�w�#{xS�o���ji<稺�?��Sm�|�"R)05\��K\-�*�pG���*���m�5}�Хm��"�N0g�֩M� ք����a�q@�`@�9�rș��x.�z�&,�XlxV64EB    1760     5b0Ɇ>�L�����k���C�9�FQg���X3
I�|,�.�wD����G�>2�E���aX�e�v�ׄdOn���z�a�k�v�s	2��$8����-�Kzo8;�y:�6��������1y�s&�O|�:x���a�MF����n,C\_��80 ��ՙOGc��-����8��f�i��f���0dW���`���fl��\h�]W�J�\�ձ�g�H��L���������ִ�)��ס��t�r
#��pѝ$툵 ��\hD�|%|^�1F�O7���l�"����J��l�1T\cF=�G`j���1��|�������ت}_�/���jt��n��F���I�F��B�Â-ݟ	x?��H&~�Cz��∡��r�&�fV�����2�iԧ�<+)B[3'��,i$I�v˶E,A���ТГ�l���q\�hl|��5��sB;v�?S}.�k����-�� a*7�nz��s�~&ҡI�\�
O�<2�j�i<ߕ�f��!b���D��j�l��V}[Sw-lf�+���͐پin ��Z�%���a�����Zi����I_��x������2#PHb������u�f �12('�+Q�����`�޵�Rѵ�W����'*7��:2/��VuBע��
.��e5�b��ڒ��9$3�ꡄ����s�(G�P��j��z�X0�nG8��z�/H��$ﯴ�����In�����Q��]�TRS���4d�C��7Oeq�Hl����c�E��O}�T�c(��W6�]pM��v�h��G�҄n�Ӂݵ��_	q�
�+���w�B��'�:���~\3\�y)l�,�FS��q�����3����Q�ެ����z3F�<�l�F��1B�iI��_����U0V(F$��$�e8�鲬ٰ_^L[��y���CD�P�܂B����ټb��3�dΑ.�oMw�6�/u��{R>-X*���T�t���[s�����20Of%�1��CB-[�o��Q�������V��������<|d7�7ͮ�� �U� �8n���zТ�/>k���f�$l8�	�I/��'/���
�:�D��`ۑ�����is�+/*�m�^'[7G��/���?�}X`k�W�Cv��z�0;Xlls���s?4��!�6�l�=PP+]n\���y�H�y�۳�ci�ɔ��"[�&���!$�͕�܎k�-��=�I��'�O;�5���T�hY�;�Ťy�JY�!����f=�_�q��YE��ϟ2���?� �;7�f��k�r�v��ϑH/�eg�]�Mߐ��о@�A�!0$(��c;Jb��Ka͋I�fp廳i��!��䏥���3T�m{��<5�-���zҒ�95?��I���= "�rӹ�`�[���3d��L2J��7f�g����� @i�t�Qf����s+�