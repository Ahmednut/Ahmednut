XlxV64EB    32c4     d40����vw�+}�v�Ig��AU��6�[���-V���t�� ��$Y>��N\LeI����¤��Jm�i3e�N��Y*� ��I=y�G5���p�L˴.�͎D�i`��c���5��XU
pv(��(Y���me�:¤fC�jZ��@1�$�x��p�6**��(�e�ϻ��1ФwF�T��@����-��&##���+{A�VP��$K���d�c�-�Ә��~;A���ɴ��J6� [r����!4��[�_z�N��<׻�J�7''1X��[Xv��$O$+�g`��G��������@џ-:�1C(Y}Y?O����ݐ1����x7I����,B�O�ƺ�\��%z'*ڳ?X'*�l�o��o]H��^�,� ^��@౅U����Ib)!vjC�.�����I�x����VI���:Uɹ_e�&�/L�J��Hl�c-�^�K_�k4���
��j�Z�e��ͬf�)4���^�e��Dq
�O������,��d�"%��8��ogE�P#=�U[aR��|�~Ч@�OԼ��kyl� R���J��֚&���5=WH�1�\��Ɯ��܁�|X�L���SQuX�6�zS��{�KU�]s�{B^��&�)z��m�@�,��y��^���0%�T��I��#�*2FO���5i�h����C����M�xf�L�#ą�����D��w$Q�I)J����N�?�L��$�gZ?"���G������c�����K|#&�96������LR �Ҥ�d�%��H�<XJ�q!ڑ��;��|B�LR8jz�a��	�O�Kmz��)k]��6����b�}bg��!\mZW��z���(ݢV`���V�U�_�+��	�N1_��&��5�i�;��,�X_(#���ڵ�������?A8�h`8l����Y��4^��M w�Z���2�:�Lg���J��	oe^r�"y�h���od���)���Gn�
��@9�~]��J�a�ZS*���5I�A�+�.Z�f��~�h��K䩠���6MI*�U�w#[����s�O>���Tغ����$B��0	�ߺ%��us5����o5 �7�2B�Q�j!����۵;آ�H!;�?��4&�LS��r#:SP�3[Z�y�G1�wtڕB>�
M4�hU�� :��h 6�/��U��u���_���a��#l������\fn�1{��tjф����M�9dW��2@*��8��L����LM��3	=`C[���:�"@��f�����������M��gh���Lނ�� �2k�l2��U���
-c"��4,?c~��-{c�	��ANw����6̀��u�F�`-�+7(	������rS�̻_�*�	�~J�19~��T+	������Kl��h)�MB/��Vj�@v/�k&!0 b��=qo�QxV���| Ҹ7?gm{�^�m��6��P�.��*ݺ�g������'�o~9=r haJ_X~V�5��8	����)j5ϼ�d��.�f���*QH����ePbr�E7���А�����%��,T�� [�⋁�8zef#���s�Z{��w���LC�8�q��ļP��-w�[�@ɔM�i_�X,��DJ�ԛ-�V�_�����讂�6x��`��|
O��u權�c}?�?qP��)�K,��
���R��w!��N�M�"�H�3���`D�{�wP�d��<���/U	r>N`���Sr&2�o�.Ą������uX��S���dR��{h�+�B��@?�DEd�p����x���%��K<<Ĉ��*�1�<��-�ɞ����=ҋzWc�)a�L;v8D�S0������Xћl�1[֒�V��2o���!F�x����ߢG�h�Q�,keh�v�\CI�1d�	�h���hg��a뱼j۽9:6�ӕ��Zi5_�e� py�#&Q���A�l�a,U���M�εY��٢���#���-CC���?�%��W썦���]�V'�د�g����G����8����.8θ��b�#��8�7��`f^_���ߌ(:_;;��`-�.�I#��yM�1s�A�o������m�M����Ώw��5٢sth�ϲa���ȿ����k��Mq@��ۛ�$U���
z%r��N�~O����C�E�V{o
��UJ��%�0Z�çXfAw�r�+�4X�Uل�<�ݐ��mJ#���m�sG�jL<��x�ҰX��{���Ή��z?X�!J��i~x���o4�<x5��h��&�����	q3���z|+�C9��J' [I�~ܸ������O�NyN�"�r�"b�0'2���P�^����nψ��_����n�&r��*f�oO���h�~�ӌ�ǐb ���t��k��h5�k��I��7x��.dT^O���	����hz��B5�L0~�h���\-l�hZ-��׮��?V��z�@jߌV����6}LC?u����C�3�"mM��Yv� ���Z-8=��O^뾼��|��^��EJ�H�WN,�x8ksۼ�j�e�T�D% �m�y�X6'MF՜�z.��kz������:.9%Kj��]�T��[~v��cӆV�oq\O�v7��æYO`ʚ<甸_l�}�nO����y����J;{o[I�e:n6��ΪW��?]�D�X��r�N����N63��_a�Jܷ�0 �XKG��Ν�+��N]�3�]��`�g�_�x�T,�G{��,�E�߲4A�F�hlH=��B@�k�ej���\�fH�eq�!q���*��B�WM�[@|�#����>�V{ A=�\'��^�.8�c��+���v�a8��A֔�J	�'�°R�^S6����ɜbb�
=�xtƮ���Y���J�L�0��w
(���玠(ٶ<�(එ u���"ڃ�r���Ym�>�
��]L�Q��^5��@	[4��}-����J���TܥI�Y�����w(KSrm:��5����C;�k�b�Ǹs�{јS�GސN�f�>R�̶���=�̊�o�97�]���q� �Y
G}<�];�U0I�fnq�&�i1E�OF�)i�m��=s�lPaJ'1�'B�5��ծ�?�1�"P>wV��R8kv��hh���9kh
�M��ɧ��2�E=��)R�c�=�M���"��6�"�G��Z=!���el����A�lծ�Z��㲾}'s牞[�?S�K�q��ϑ�VL�	���T2�U����M+ޗ���6x )�+�Sx��ׯf���Z�FBkv10V�>��33DoG&["z�Ax�}gD/!Qz�3,)7C�Z7��MɣDf/�B;Փ �ĩ�Ne�)��.�[W��$ٞ�w�;P[/A}�n�