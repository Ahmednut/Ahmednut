XlxV64EB    1e37     a80RA�H���jF�9�Ih�*Q�m׋]��=�<���RL�ej'Ҭƥ� (����rcdM��KY �j�f�]/5����2��48]GL��ϙ˕ulFv��wmq3 ׄ:+י�����r���B��6T���E�G���AέY�f�yB�Q�� ��{��A��?�S*�i@�h�ş�ea�� *R�;�4��[��o)���R��?�+~yI������js��
���5�d[4Kc�"%~ۭ�4o����9nc��/��F�������c"���-TnxRar�O���]B���R�.����=3�ofs;QcOt�a�?ãL���L,t/�dr֥�"�~��
�}��7�e;g�x�OR�e8�c HL�f��I+�i�,��.NfTv�I,bn(h7���@�n��|?��x9Xmء������DXtWۏ�P���R^ZTu��C`{h�ٌ�����7,���/+�����MIQ7���U����)�.���s�<9��m.��E��F��'6ul+�S��rs8@N���,$��)�^�N.ݶJ��gK��"R�BC��9u"���T�)[��<�k̆W��\�o49���ky28��ri�%N됬��jr�9�A�Q ?�O�~Y�����f���Z�N��5{������mv�8�.t�x}��`�ĭ@`��No���ይ�Y�rZ]��+:��N}Z�ɳj����s�ܷ�V�gs -��`u���%G4��g���=$}-e1+O�@�f�&�
@�Jʰ�]}��.?�0>O���j�?�h�o����`$�"�똟kh�?�,�F,1������k)<���AdO}p�TEU�_٣,K� $f�\Bk@�,5�5�zQ>_�V9T߭���f�Yn��ch��ڭ��<������3�O4���لT�*�v%H�>eTuC��6�c��L���R5�Z�}��ŒL4̼@wL°�yKѶ2'�18�iL����6���53�D�m�p
�$<3Qسx2,jC���ZPR���Q�&��TcWf¤�[�Y�¬��Y�c���N/�͖C{Z��2}����R^c���S7C!�Kb�PA�"TB*�����;#ǡ�!�=�<���O�,���������_-�o�R�G�qK|��
��d�.FW���a
���,~!V�I���dK��Q�M�5\���:D�)8lY�\��g����[��psRO)T�Lo�Mz�i|�{�.,���a�4�p<�TJ���K���{I��Xe���ջ��^�Tq���$��8
�`�=YF�i0��*�B��q�G]����7��ty���Wv�ı�O�ds0��E�K�uZzԏ�P���Q(�?�`S�#�vg�(�^�'
k����p/TUR[.g���b2ԈOHajl�<k�^�v�m4:�3!R��&�8�rz%��	|5�3���$���ۜ���Q)�����&;�#]\���Z�5g��Mn�mj]����Z��j�ƭX���n0�W�J,>�?���q�U�.�^�L_Т�w�=_cէ�(9%�s��H�&+$^��ز�*m��ykeg�gBs[(��=*NE��U<	��P��Of6`��qt�Ѿ�%u9�K�C��O��"UuQ�0v��*
]���D�O#��7G�d���ƾa�0D�ɬ>��f��l��{pv�w�!'�e\�K���ф1��Ɉ��؜/Ml�/�GR�x
�Q���<�jv� ��᭦=poyK��0~��6.���3U��ns\:�����8�y�Pf�A�C>�M�@��!;곪p+���SI2�5�'Cl^��8����@�R��[`�m%��X����!@��e\\�<}���g��?�X$r����"T�<5i~���_�������vQ�6�!}���/�����.�*_�� P��L�ځ�����+�ԝ��g^[k	BZ�!,�L�����y�r�	qD2�YyD����(5<)̦ =#�F�PN� z�g���j7ODI�e"�i���U.J5���{�b._�N@��K�ӡ! �N��x��V��7�#_Dl`�ؖQ_�~�]��,l-y���{8�P_�~8#�/��ߏ(��D���w疕��&x�l/���U�&z��Lu����'���:�W��S�Q�Qp�u�M3mo�+ڙ��U �����̨ә:t�`�N�Hz�����&�P~�q��
%Xt8�"1��r�(s������XIU�!w�U�a}x�,8��/���7n+�6E�ɞZ�Íqxz�r>�.�����#-� b�'��մ	��W"�s��R�����1މ�- ��gU�J5�{C~�h�i8k�M&�M�)ʙ,c~�"�x(���D��3k�f��\���&CӖ�nH�W�j$�f���}�~�wUk2��1tO��%������m�#8�/�l��E�ߡmķ�@�|'�3�&��]�H�4��;��'<���Y��T|I����v���~H�/0z��fH�N������j������B)Lp�[���HB߬��ww�0i\R��Qv=�sq�>h�k���sY(L���A(�L7�h��e@F��w�WE�g=y�q� JK!�J_u���Kp�l[�\L�Iӻu��w~i�4��G���g�مH��05���x���k�m��