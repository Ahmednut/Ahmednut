XlxV64EB    fa00    22c0���W�GTU�����'�V��.���GQ�Z��g1K�[��rcf'5{�����\
� ���u�L�(�`�W����L�\�X����d��,��CG���g���*a��������|i@�U�L��A%�mt�tx�u�C��Zl�tS�98�uI<?�����~#N�6P�����	(�]�p��*t��q4�c�bgC���ٛ2a��Vy��'~��쮠�/H��.+�	M�Y�����%��:�g"�..��+�K��ԻBԵ"��[���;�d|��Jk�!ϾNjd�$Fo�]13�V38�r,�׭G\
"��G���j�g�GH��Ua���А���^�c�5?O���-$�F�2BNZŨ%2��/�*c#]���[g�B������R��^�J��&U[#:�� �3vT0K��Ȼ�\:$+[�-�����g�� ҞF��4��q� ��&��Z�ЮI�$�����r/�& ���;�4���Y��8:QӇg�SKt����ٿ�'A��qI���-1��4��
koa[l�To 	5���:_�)*���<K����2vI��?5ՙ6�S����}����	��+6؆Ka�
��Ưj ��$�*��}T�T�D���l�uV١��K���!Z����b×n�^N��g���N���3����1�B;����kw��x��װZ�{�1R���p�^��qI�W�ɝ�(tp�ߤ��Z((cv��x���\���5�ܹV�)�6]��/����ؓ�uT���w��-�����o(,�`Z��6��/I,�F�1> ���E�a@���a�) B^
� ��3�|��X��'ǂ�T���;9��W]����-�e�<����F �Eh(�T�BH��!.��6#D���d�-ay����XnRuI]ys�K8��Z������M�i>�0Z� �^��qi��C�eHA��}��[�(D$��ޕ�0�\�[����7^���8�ʻVY�~�B�`�vB��"�)a�-hPg_�((W���U͙N>�C�I�\���[rO���x�x��>�W	::�-}6�߽C@#1Z���z�9c�`��O�2�
���wn���JD\p�X�<��~�"{w�Hf|[V*�'B7���*h!䇕�ϖ��^��t��w��7{�\����4�#�Q`h��z~�{&��������`S�n��y��fT�D0|���&M��=��mUw�3���Aʠ�sA&{��q:��hگ���~��4�M� �����@|��kϢ��/`�i�}��i�=�f�P�.H�=�T"��_�U?�����d˵�WϢ�6�F�^�-�������J�В��K:e�L2;0���'�xMl��Dq f��^�[�֝�u'H�D�h�u|��hP���-#A(LS!�j�C���f�NR�t"��~��k]W��J_@Q�H�a�8 K��Ì"�������Adۏ`�0&t��"��?�}�/�w7�� �A���=ͩ�E -1��8���z#���q?-C�#�o3�c�5���ĈhJLm����F05
��YDnǗ�$�޵P��fer��-p�G�03��s����^�S͠�Hĩs��^����8o���Yī§ƣ��V��fsV���cT�����;?��[e���߹��/|�ã�����I�~8>�~�#�g�����`0�$��$��m�0�Y��m���F6U�C*>��i��FU�M��+j��l�s�&�q�_���~9�c/D�ױb.�b���)#��)?%�AL�G�ϕ�	b�X��H��
}�c*���AOfe�߅jbtn��rmz�A=bط+�P�ӛ�V�qFoCϢ�9�O%\!B��������e��yw���K�% ���X�T����-�V�q����	��Ԣ0����-/R!L�E,M@��^]vˮ��),���%��C���fKH����O���RP�n"��2zh�%�O��>����(�|�e�|����Z�D���J��w�Q��I}9��Ap�c�b�|��jQ�gu֬aVx�4k!�鉇Ke��歆C�	uU���F��� ޘv�lQq�Y�pѱ7xП�������_��p6�Ֆ�m6,��z��6
�cJ���O�����.�2婒_f��^�w�=��1��v/�m����3}��h���M��mb���{�ۻ�!p�R-0l6��je�r�����i�KO���%���jɴ�ϒ��N~3�V)��n52�s�I�o���L��j���6�i�n��d�v��K�E�	>
paD����7+����ȆvjP4�Ɩ�豀7 �&{hW;�8��.�˪��������W$VŢvz�my/A�D�����+�0�h�mq~��]�0ό���a��2x�ر�	�pU�~���S�ω���w�f�o9Vd7�V�NR�����P���ͭ���"~�m�$n�	E�=�Ӭ��9!;�U�ќ�1�29sv����[?���Q��#���^��\4�]��+aPcOִ/�nc���p2|Pm��	~�i�*\
*�Z�"�8?�|�
t21�����N'�rRN�����%�!��,S������mL�o���I,��G3 l���_���
�8��Z2���i�UBU�Kao�a�^�a�g�H�,<�/�Xv5\C�M����e3FMܼ�(#�&r��0=@(1�wr�����O�m"�C*5Cꐎ7�n�`�M�s�Z��ԩ��VIصF�����if&���8��Ө/X��4�wκ�4�m,��{v`�0�f�4��DQ�tri��=>@}u\��3	�>�6Z��[힑*[�0��vVX�B�G^�9�~� ��O���ҹk�� u���3eY�b,�Z?"�7v��ނ��W�EC^�f��o�5���)-O��K6���5O�t��9��M���#4}�����sЎ�?F�������'�O�������#E��|T��"Us� �}�5��7�	z����"G�U� z�Q���c���-Z���s2ˣ+��w�~�'�Gg��u<r�[0D�1j:\\3m��N՜���) w�J��ܳkg ��Y�1�-�2��lTM�U�MB��U�M�� �ڡ�U�ӣp���۫��EQ槜����Et�X�<<
nEI�k'<ɣ/-3ZL�x�*)�����i��Eԯ^|r8P�fD/o�#d-s��r�^�д7��&��cq!�#�]�~dQ{� �\m�ᚁ�x��׼,��~��
��Ը�	~5=8���6�����G��R�����ݧ�8�wC8r��a���{�B��H1��I�^������� ����ْ1B�	\��>;��ҭ�8��(�� y�L�CA����3LUX��$��r��I��@zۼ�]*�(���:e�����{��6�P�eʏCJu����
����Fw�M�RzlZ�gh ��f�g�WuOj��ߋ7a9�'R��d�����u�6>�fO���D��f�f��1������k��u��h���'�i�ǐ*rsLD7�<-�����<?BO��2a="���NB��	{�TW~kMh<@�gl#�o���+�}ᦏ�s�;��2�q>���]DR&�5	X�d�����d}3�Թ].�9d��K��hد� cg���F�jzO�~�b�a�Xp�L]���]!�W�� ���A	kWnW�Ro���$�dy�����gVh��5EU�H���|o���Z��t�c��K��uA�"�U�u���lQ��,������DL�4>��f���OԀ�2�Cǡb�iN��C�C(������%S���Ӥz]��M��;���wl�������^�n�?�82
]�D(3Q�p�������0�h�ix	��-;�Ԋ��r�vP� \U��܏?~�x�}L*��l�a\����;��Lx�}zЄ������G��a�Rim����
����E䄝$^��Rd$*a��*�(Vo�N �`���F���o�@��Uf�pVw2���E��`?V��, ݼ;u!3����(mK|w	n9E}f���qycj�Z-4��U]�U8L�N�kȠ�hL���2�c_7��C����L`d�u�� ��-3�LF�0T��r��U:.�2��H��,��}�\:\>򭠬I�Ι���p܅*�,
u:%g�D��� okwC�=��8�1�Bq��o�������]q�N1BhB�58�}�H�r�B-�s/��u��:��C�;�t�':��C���ս���E�5�o���M��)���Z�c<�ͦ�$��̈de>P2�C���_0��ߌG�c-�5�O��Yw}�@�M��W�B�uh(.(�Uik�B�mbeKvݷ�̤�v^n]A�6D����W�
��h�{
7#Q>ߥ�v�6�
v7���Қ(V�eGׅ��X��}�{�D�*���[<^ǟ�_��zaC��Ƕ�KJ�������ؙ��Sw�����~��0q.����А�������t�,���_ׂC�I�0�-���dywsɭQ���6q)�.�aZ8���B��gߣ�?;P}�������+4��t�w�,�Ϩ�ӶTv�A`Ǖ�<�N���i�[ǹ[��Qz�j�>����$�x	x��ħ��XZT�z��(��1Д}2�U�m�y8BeAN(�{)�C��R���CI74{}���7��v 5�w���AM6��xfhZ�^��(/�����'��g�<�'��v|�C��OH6��;��yZ3���i=\��6��t�J���á�&`g�-�;Dzf�ӅU�q;e��>�����
���A1��5;��Q�sL�:`UJ}�r� )Q��yD*�U�;]UXP�p��D�cT���K����<?��e�Ì퓍�^.�Pk��&�a��(u���S\H!�5���:���[�3|����"�`K��~��j[��b��aɢ?uV���銇�&�$�$ʏzRz�J�ĸ^eټmX�97���2��k����Ԃ��d��eiBk��{��#]=.�X��}a�}�*��!�"�#�3��B���ׯ����i���G�|Z�Ƚ����� ���@U������w�V��t2%(g�!��4ӬCF(;��n��l	�)�&�|sca}��%E�̒����.�ر�Q���}�f��}:�G����*y��^(�r�w���&_<��Ⱥ"-�*On�k�'�=����/|�v?(j:B��ׅ#SoH�1{��x|�z��-9���Y�}zN��.a��z��u�&g������%��+��cF ���(g��F pEm�3�Ԛ~�\H|Rp�h9����h����[G�c-2���y2`����_+��񠑞��<�;��X][��:zv��di�z�fFP;d�@�ng�x螗0 
j�P�����O*���[.mˎ���w��
�ɂs"C��
L�]V��6��C��e��_?LBzyg8���3XI�I�#M�������yp�C5�� �L�B�".�.{�2-�rQ������	0|�;}t���R��	�9#U)��9��r�ހ��w�R�zb����F����T�e��HuO`����?>���)�B(2a���Fw:��kv^1���2f2*n^ߘ�Թ��"Pp1xw�漚l4�2�;�I�K�f�1�]�8��=z�UX��a�¾٭z�������[*G�A�Hً{l��=�e�������9�ٞ�p�<4������S���Wp��ʙO�`��8�6e6�2�,_}�H-T@��6�䊱�T�"�Q��~f��Ո�D(8�D���K�֕fJ~��>l������*��{&J���Lr��I�Gv������ĕ�G�۔7��^���~�8;�����#ᖵR��[:	yw�+E���XQc��Urf���&��L�zWO�9�U�
�>����xF��_Ɍ�Ӗ��>��8TH �x�F#�>��*�����/Pa��1����Rs��S0��D�m�4�b܌�>�*5�?���~�η������Uٝ��m-fsɯ�Y�1��s���r�s�Ȩ�݁Y�+�=`z���w���哈�-��y�O�wl�Q�(~�􊫈�s�! �h��nJ98&|K���1 ]~�L �b�� :A`�h�H����3��<}��7<��6��	u~ۨ�%�����ȭ�T�SNz��x^-ro/��d�k\�X��`��|�]��1Ы���3E�Ԁ���ѷ���ܜM�]] w�`L9~�K<n�ϮX# ;[�I&�v��'&������G&�9�^)��ݦj4�993{� ��>����_Y��'��Ex��l�����B������e/(���{[0B�6?yzE8���RD������@{(Ġ�M�$ȯ�>���6�w�����xvу�,�#�au�b8���'e��DHź�?�fBA��1,��!҃V8�~����"�X��Z�U��ȁ�^t4R�8�o��<����.�Es���W�1~����A����'����-���m���q����V��tu"u����d�3t�ӷ`ԑ�4@���i�;�4�NݔH�f�{�ĂӐH9��8�C��ZtAs�3�#L�|�tso��PqO�1.��Qf���T*�8�0l�
/.^[!!zR��D�G�*C�f��Y�2��|�)n�b{_og�Om"P���������hE:.o#��p�������*o.�����z�r�z郎+$�Mۇ�R9sj��_�P @����=K_�K��r�݊W�H����(���EWh%��	1c��7�~Oґ
`���^�dJ��uA��	�.��N��1\r�8��1x.��C����a�L�2�_.�h�)��[��Pi��=�3���h�f���Pv�_w�0�, ����7�S�ꎣ�����X�ǽ�I��2����"\#3��f+9X�>s��쁗3{�3%kl�-�g�V�Z���/��M�����x��=z�_<�ѩ�����j%�%8΍��������X�O	X��;���/�CXXn^�ݕf��{+��V��i�Ml�#���[(�Rޣٞ�{��Òy���
�g�SC���JZ�@��p�C�zd3�R��M4�Co0� k�H(��Ѷ�"[���y���;�V�r���:/��`�(�$�vDфF,�tm�O��v�"��³9�+�)����vu���u�m�@��{����	q��L��>�A[�=�n�S�Ƭ����W��:�xlFa��M���M��N��mf�	�U�
`eN~o�������?��շ����+�ͣ{��"��].WJ�L7ge�.{8:ulZ"��5{%:=zL&�㽻�:n�ŭ��a��!��#
�<n��I���J��Fb�v��V��,�[�NS���5��oV�U
�a}_�v�<�#l�
ΐ�Y����-.�[T��L�/.�+*ַI_�}p�������	~�w�dﺿ���XՈ�u��ծdr�c�12ZH>��{0�Kb+��[_�#�Ⱥ>���>���a��C\�M���3� �5|�W��R%Sp)O��H�����G���M�{o� ���{wG�L���ʽ)�B��������p#�e�3�!��f*n��C���� 2�X묨&�����!�ΠF�M���/,L��!����DE�(raN��E:0�nл�w�ɛ���0T����H�A���w��8������pN[���5ˣ�S�u]#2j�,e�3"HݒN���F%��p�˯?���Q��8�w��K��zx��W�{f 	�'�.��y��Kݮ�%�)�Mr'lv�`��KmѦb��O'ή|zt24R��b�b������0U7d��~,@��A��{'�X,^�`��"!,K�#rƈzr�dF�	ޜ���X<V"ᤒo�_E�#��y>4G��|7�9#k��8��R������vH���=
�$�������jB��Zy��Q���V̫�H�0׈�D��v�I�e�#���aZ���-۫�z��� �Hv���b)��;�ˋ�%�q�VU��x+Uy�aI�x�F̡�C���h'�E�4��Ȧ�U|h���ڍU--�al#:o����)wR�_�+���$<�^���r/�G�JA!��2ռ��"&2`��=�}��3��0�	�H�Pv-�hS�t�FTz�� �M0ɥ`_o�**�p�P\RGO�K�q�Qo����&����������'��d���9-Rl�ģX���*s<���$8|q�Iw�,�N�X�KL�ܸ�<�L�7p+ԋn�{�^�yH��&4�zʭ�����toV�p�}[�������7�=��l��O&}N[��!��\b�$�:1��Ua��/~U�ż�&Fxm9Ľ�I��C����/�?3><�x�z#e�ph�K.1,h츜�O�}�Ex����Jh0b��L�N�̈|�'����}����C�M+�3l��G�Kܴ�H@��������j�t>�]X슀&a�",R���SHŹ� �b����dT���C
��̡ve�[�4C��fON���4^gV2k�	��Г�l��J���8�!���e`���	O�J��xB��V��������9C�W�j70��� �
~[^K��uz�nt�^�9�mK��%��ӹ�d7����p@!�%�r� �#��x����{��]Ғ�b[+�����b�X��mM*��9L�
����ʖo)���i����8a�[�����J���j����KXlxV64EB    fa00    2440X��+6�ў4�O��!�nE��O���b�U�8i	d�"3h���
�Mf��Q����T�-���8ݑ�{}�R@���U��v"B�]��Q��{�*Y�[u�c��-ƬƜ껖�D�l�>T�rg��ߣ�|�fq ��K�0�.��ܒNxN3�H�5��B���*�ƃ5�q՛��8�)�s���J�r�v�ٗ)����gW�9�����uZAh �����{SТZ��a W�k%B1CMӳ�!��ȃz�#����E\�8�'�����X�����HU!}��0j�3YTx����g���%�b
k�q'`���_J"#��e����S�'Gn��T��5��c����9n���)2��' �&h* ��	��+��;Ŵ�6��_ G�� �*�	4wҡ�t��QY�xk=�M�=;`:�:� e��1h�M�h^��5��w�<��yr�Zj?�	��-B�|�X]v]BJ�o�X������f����&8K�.2���e�X�!Q�d�{[��-�t��
����\��OO�HKם�'Q�r��K�&}��-�RG�:CW\!Q��fl((����������P��V��ǚ��@���_�t��{��4C��:�OYj������T���ڬ6LX7��*[@�/Z_�QqeL���F���C8z���b4��m�5��᭾? ��=�5����E ƚ��*��Z�0H���,�0>[YbU�m�DΜ�H�2�q�a�9��uf��I��1�WR��yȬ���l%����m� �� ��|@�nԱ��Ƽ�D�y(��d
�-s�*�l�_G�Z )øp'�K���g@�t$M�4�[�~s���
'y��m��9�T�<olG]c���t���N3e�����"N"EU�C������:�%�Y1j}j�㿖���,=�.0I�ݴ(�}��:�W����G$g���ܝb����d,�Q�0��@�N�O7����M��M�����G�n"\b��-���$����|`�t�k-�݀��Ij1gV��E�up�a���='�^��1'g_V[�c�M�I-���#b���Bǹ��[&[;�3�:ޡ|dK��S��	'_���s.V���]�=q�dj�n0���R��'���ɡ�����^�xjg[��署E�A��B�<�\/v�*y��npe(��o�윔�;����6��\l)���"��.���b����)�HT�>?�L�ː�Oo��;�H �?�.ȁ�m�e R<�>1��C�$ڿ�%gy���	��G�6�+��v5�8A� �#c���:�3K!�T)?r�K��u��,�0��&���u��S"ٚQ\{"&�;�+�"�ǰ㨃b���}I���A��*�W�*�B�#Go���L���X���_�/1mCo���=7YͼiE�+pOTܯxY7�tG+f h>4�˫���_�X����'N����T�j���y{4P�,fz^��G�R��h�t?����_uvy�7��.Yy��>�J̳��7.���o�?�v�t�,�j9�pxz���!$@bU��s���K�d���,%��U��{?'��8�2m@�PjQ�{���d�˨�`�[��3�;̓|7G�3"�`YC�A������,3we)�wA�<B�e�I���
��Gě*ל>u�<⩀R0��^��۵<A���xm������<�@!I�5�t��D�^1'��T!��^*�НJ�-bK�W�t����$��vg�f��X	�Eh#t�<��v��
����B��7��d;?�u���\�b�xA��X}�BPW�l�y����p8m�,�?ǘGD�Ӈ#,yH���Ư�%�d�rW���Wo�yg��B��7_�ؔ
��Ԥ��dj��Hh�ؠu��sm�Z�G3��2�{��Y��?��^!����=���}ޱܨ�=�T�pg$]��d��!��q�����]���*�t�m���n���nW�f���Vz��x�	�'���Q���I�C|f�Rg+k�:��-}m��ؚi�ˁ���sR�Ĕ^���5�T.�p�ʕ���<A�������1\ w���s����^��%_�х��Ey�����(`���j�;�WZ&g����iQZ(���ǫt4�F�d̷�F��x.ɗ��b���EU����C�F��
�Kgз������r�QUP������ѣ(��e�5ZG^7��L�o�F�5Θ�c䕓�<K$%V�C�Μ��+w�P���v���z�#�!h�0B��gKu�q�@h����$JfY��C�����D�5�lL�R"�a�m1E�
&h?f]4������ ��H�� �	8�C���@E�L�Sn�w:��Ix �*�c�^4�}�-16��k� P�5O�M����;��*s,��)�ӻ�C���}��mH�{(�L2�X9�K~�Ɠ z����
e��hx�+M�����l�� {Y@��q��]L�"Z:��~��s��8���?���T ��`ؾe�*�݃��[CR���}����8�ܙ@[<�S�&�u��ݖ.V�+\�M�;׿���R֖��i�?I�;�	�װ����9���K����-e�^��0a�$1���rx��/u��A�i\��^Ѓ�_>�.נ�ˤZ�f�V�3Hު���~�6r.��[�:]��Yb#�g �2���i�r]���X�׮9JY�����Z�;�ҿ�*Up�1�-#��~�BY�Z�n��ƿ�T~UVd����/[L�;�
S�<֎'�<1�e����Jp]���=��!�gS��r��>���T�+��2�;5>ƕNX�"��<���?�r��=$�p'n�p$�\��z�&����O�j&�^�շu'�r�8� D���I($H��;_+|lYr36�ѫ��3��-���i�A�iT��^�w�x��E�(N�,s��E7�(/���ټzJ}^�r ���X�_��q\O";�QC(��~J�p���q7P� �6���ZK���|`e�_ɼ������/=���C���hn{���8h{�~�7D�84:+?�b��Bb�X�
�������v��>�o�[d\H�T�?�v��!����TV� ��K;�E����JG8	񅝮">�� ۇ�1�7�?�
�<r�"�3L�i��;k&X)��Ҙ�6z�R&���w�Ґ��Q�Y�!�� �y��nj�,c�8�:�'�����I�F����P�>�ݜ����꿟���D}?dJhƃS��PĴ����N?>��O8�n���9z�qjT���U�ꔿǏ��n�HfG�Uwў�Q�g]q�l�����̩�s���pʿ�2YCx��j�%)4+�܆p��	%-��b <�k��:j�'�g=ą��Z�������R�q�@j�gZ�߃�sl��{"�c�"qSg���8�>��U�nJ���Pr�<A���R'��9N�IƲi��,=^������K	�=*_u%q8M{㲶>)$z�..ƍz�HY�(g��6���[v�w|�`l�60�ګ�pC.���G�e��	Y�@	��4$+�DF�q�@M�� (�T�LC\���j��M�W!
uu�!M�p�kr�t��5����#:7>��<�����?�L��qv瑹�2E��	;�Wп��F��>_�������CcKr�#�{��=��j�8��^�.�U󉇈�{."?�H��(r�+=z[�K���;��-���k�1t��w�_��H�� �U(�=��z�_�����DH�N\L�N��K��NDP�1�%�k�Ƕ0�+�QR�ABU&\�㫮�VVf/	�I��3�V�iED���ݡxz������|�5����<��Z�xotsکn���wm�����TEn����hc	�J�p��3:@J4�ͦQ�}S�镜�Zqp��!���1~_6��%I߱:�jّ��U����7H���b;cM�~�o���?ҹ��	n�G���VA\����=��\���\��X��Cn ?�;�?������A�� �a��-_N28��
��^�Z�<���âB�;9J�`󻤘�ψ��/F��z�U;$W�˽()+�aM����y�
���I�o��&���{�e䝺��CؔI�zfS��_A��}i�]�����Oy8j�Ԧ:���-Y�ƾ��9)�,�����t|:d��{�vp�x@�J��djm�A���|����|�g|�f�|�ۤ��=�3���g{�̲A����]	��w� 3�ğ#��EE]���-\�E���ԖA.�V<<LfE�Ób�]��=��&_ɇJ��ꓑb=�b%��\�/��5�E6�q]�6������9 �7L��e�dX�;�\ĕ�u%۩B��Qo���;Ϝz'��\O�<��:�֮�3�}oWc���K?du[u��A��*=~b�Y��8�V�[=ys�'[A��%�__s��aȀf-�����d�غ��k�!W��G6e�tr�gܯ�m2����(���1N�S̑_�� f��2���E7�f�'�dq*��~����;	m;�l�w���飗�N��G��kjQF]'����lG�V�̽��~ �z���ޅ{,��Y-����MH`Y������ِ����i�-+��hd�z��%��:�B�q0�w�W���W.���VR���E�g.n�r�*&�L��f�@��������N�H�s;dQ)��T�y/��!��we�_��'�P�땾 3�ğ��~f�̂/F�_���ϧ"�1|,{T��)��/a�x�]�P��8����M���I�_<4U�Z/`k��Pܕ,���<����Wvz�U�x�����f�g���� ���/���:T:dE��4��°�t�5�d��2�N������p�I��S��^.���\�ygjAW��q��Z+|7�~bz�J��%��v5s�B���Au��d]+r˥��;9M.#�u.�l}#t�V�3؈|#�K��,�$��U�/�J�gJl�h1�v�����l�����G*��@���N��A.��R�2� '��=b���U��iN'˔�fz�����G8�c��>�,��`E?���{�Y�H�e
���x�b���,��k��#����"�o)���_���W~��!��FG�HS>R�|#ı��VP��x�y���{���I�r0��6��_G����&u���`��'Չ�^5�j��[�h�,0�^@/^J8	`��s1#o�� ���O=w���$A����xk�%�j) \���6H��^���MF��(�,Y��}�I،ij�������s��w�m�$��!=�G����A\�'�]攉�~RT�����6����}U��iP�?ص;��XotX��_3����[�`�b3����B�spB�6E�6��oe��"Ǖ��Iۦ��,��$�r�OΘ}�D~�����8���t�P��)�E���	�!T�EӸ����ؾ��`����Ġ�C��u"�����Ϗ��m���ԓ�Ӫ�t>�O��+�qD�hƠ�'Z[��>�	e󱵀������|�$/sa����3��̅��u_�[A6��~W�K�V�+/��*����{`�y�*����yۯ�P-���s�S�P1�jx��c����2��1�}�g^{�_<3������'50�߲��PL���u�QJ�g�=�Q���y~A�F4�&:E^,�'RQ�>�n��#�R,v��e�g�K�ئ҉�T7f<Y�{��\+(q�˗�%:$y����x��/�_iV��A��i���P�K�x��s�	s���>���sC�n���&u�Ϥ�;#0v���ppv:�\���{�[;�F�$��LqA�׊eA�}���߻́�]�h<�	N8��
�p��`/���Y��wn��W[h˓�,%�G�j_�~�
x��l�N�y���ᨇD��W���u��t#�F�%� �J�ۡ�7dL����%�d�����I�o^��Ѹv�A��:����X�f;�f�i���8�+�p����l��6�y�.�r]�r~���X��xH�}Ci@�u	v5���>�0�}z.�.��-P�z޵�5=�=Q�{�6}�!1VJ�xx0��O��c�ӒYe�!�3��� c�2���~3�K��+n�		u�&��ֲ���k�+�4`GWVAdQ�>��U���9G *M1f�F��@��1��_!������/�i]��T���5p3�,���N�?��N�_xEe����t��fjv�����)�!��w�݁��r��r�Q�{&�a�rs�ʡ��)������B�@��ן��Ό:V�`�NJ�畏��zO#Uw"g.W��撈���c�zӎ-"܇}��xC�\?rj���r�<�5��@�`�_�E{w����&U�b��ٿYʖ�Md7/�bц�����\!l5N�WK�Q�q��?(`�?���߁�U��#�nQ������z�ĝ�����z�'���ZQ�~���y!4��������%�7'mx��XB�q^&�]�>���WGV�me���e6�Ȕk[w��}���X��{�h1��暦J������]S��K>!4jߧ!K�wV�Rͤ}u�9�!a|�p�c���SI���b.�!�����nn��c�jY�<�S���x2���e�����!r+���)J@N�w�I}^-�"�-�����؝*�*l� �r��]C�!�NeP�	��*��i��F��m��f���&	����u"�cZxu�t�_B}�Z< �;�B�Ė�:�����O�R�	�+APCˋ������"����[���C����T"�SU���,��
�R�*5�!̿�����E�(�U�l�&�[r��%�p��X�[�̼���;�OB�WsE������G��� �u���Tp1IHQ-�<?�D��M7����%��>@�I}!C�
�q8�Y� �-�ɵ�MKX����F{����Z�	�ʀ��`���b:�* ��U�f�!d�Y�&��:�ðo|�E�n��_����Ep(��d��*�c0874z�yl��x;�������A�C�g����]�8S��h�D�� �c7�ѯ\6�+'�eUFMu�&9Qڰ��bGIi���ƫ�d/�+�U�/��V��׈�I˳$�!��y(�R�V=4�+�,����n֯�%��}��9y`A�]�wu�8����g�v�\t���~����8�9C亸qr )�x4_/f�6�6#���/k0t���9<3�_��rp&��$�r:�+���� zx.�9�.�8v;�a�׈�x|�`��X�/f���Y�Ea�91��ՙ���jľλ�(��������vp�g�0�^�#x�/4<���(�l����eK�å�,W�����uT��@� �����gN����&��.�5H�6�U����T����J�3+�0�4\��E���.������-;��/��AL������m��m������-��#��/))lL��Ǐɛo�bI˾B_���&4��� ZҶ�Q˂��t������B�b������N~GApp{x[�o�B��2�M��� �]Xz�|e��k2�E�*��=��yH��nR�Ȝ�����1Or��B��N=���}9f���b����!o��ӵ�q�]gSD���WW.:`oᲵHD� n��Z�^��@�� 8�}���tX�������`4M�J�,�\7��k��u��z������~�Uz�<����}��d�E���dB	�jQ�9Z�}ݚU��09J�SJ=a�)낔0E~�N�W���9�o8��uYL�p��%Wi��y;��S2�[�kp|�hɻ0�ո��a����72ɧcv��`�������E�Y�T�3K^��x�Z
:�Z������x�އ�o��H ���Y]Z�l���G<��3 ..؛8�$�+���a�=�9�}4`������R-R���1 �}UԈ�������c�>�N�m/~��JyP�f)�^4:;1��P����5 ����Vc''G뽭Իu�"�Ag��@�t�no����j�>NNc崜C0AG:�uP�ض7̀Uڜ��v6�����dmL����o����8u,v�^ ��1�[�S����E�x�+�ӢR���σ�,q⤎n��R���LGYI>���]�b�����潘�:�3������1��C�G�h�A��0��:��$H��NdӁr���uf�cwWD�U�}rU�wgZ`w�M [�(u�Syjn�}h��%�H-��P��n>������B��M����+5>�}2�*��ެ<��G��4~64��a�z��&ި����b;�@ol���ܾ>�&
�+2W�����ǛR�q�y�I�.E�2��:�85H���ԟ�cv�}�e����EE�y��O������p��kP1�.�K5J�#��}Y�Z�y �FKjWԗ�����F9��f�_e�<��deOBoX
�}��Z��g�g�D��1�=*!{el�����;�Ɇ�d;�B�5�^-;-۳ڪ�ik���>&S��۾ǋ��%�O+�h+��V��7�j��#6Z��x�D��b}�=Ab@�)�<�F5C&������W��k�o,>�&>�|��Q^聰�:��ϔzHOX�i��J|�{Uｶ�&��։�I�w�4���ؘ)�F�8���W��l��8�}��?��m|��9P[M*��sJ^�:t�U�P���~wpj;w�JqDj/xhy3�bm"�*\a��
��Y��'�Mſ�a\��e�D0��z�<��24����'�ۧ�VX�S�(1 �
F^Op#b�Pj<�yO"����#�T�k���(Rb�V�>�{���"�Y1j�e)CK�t��ۊ�YJ�.�^}��jYR{��n�ֿ�,k�3�=����r!��YAM%9����E�б�Ts�9���ɒ�|=�L2���� �b(?f����I��z�T$�h�<�L�/�1���@�vm���N)�_�(��Ĝ�İ�a��S�Y����K�Gw�r���V�N���ae�Q��501������D�֧Á}lD��6�u��ڋ�.�xz}��Gt�5zƮg]#d(-�<��8��Ո͖�7�B��ҷ���.�Y�5�Aj XlxV64EB    fa00    2100/�=��31pcEzS�5$Op4�%���$a����ό���+��i���G��B�CT{���߷�@����T3����q�y������
�f�gG��:��pi#}��} B���� h�����2c�ݒ�a�"��� x���P�v ��z<��#
��4?3�Ȏز ���";R*�d|��* ��v�bǶ�	�L��"j%�����k�����҆�H]~��A�`��/A�#J���eh	(K��DKÆ|V�s���j�lRQf?q��>k�3���/����m�ciY|���g ���	��(�J�j��)�AWi�s�n��l�*��߈�<6���#	��!S1��ʢ��X��WX���M3������.�������%�@��j�����^K��zݘ\�̿,��4Ő��Ȩ�U�d���������.sW@NbթW8����|+�ʖ��U.�k��?�G���q����G+-PBO"��sW ���Ҿ�N�e�m��)M}�Ŭ���\���UX�mD
�qVܶ'f}��U&'	��@��Y�"#��Ra/���2���5>7(�*��f9�t����F$��qhT�I"��=�������~ ��rw!�
�c��*7[� (e�7���[J�WǬ�TFe�cj�7��A���+7�:��)v�ξ�a��ߵd%�e�ld�a
�*f8ެ�n��.Y���Pkct�_��N����_$������^g7���paR��͊N�4��c��c���+���D��"�M�h�s�x'?fc��uZ��o8��i�nD��dן�tU��\��Ǥ��`��<g��POX��H�!j{��{��R�1uRN?̱�"*�r8�\��7r�זL�,���`��Ը�۬��|3T��ٴ|�6v/Y&��(��+J��pG��Q��;cAY�Ob~�C����+T�҉���՟G���YT�Y!��N�`��~��z����������`YE�}*h~��u��
p'�F�g$ǜ��"�4�x�{�&�<��p�^j
V?ԫ���&�\�j�����y��4����_��4����3��(�8�ˈ�I�ʁ(2E��'�fް1��<��b�g�.������>�[}������޿R���ƎUۡY��1�����h\�Gk �����E�S������	��P�W8�|���[Ej�a�D��"(���^��C494ن���8���ӻE0"����rZ��?,گ)MVn��}�FǪ�����7�Z¬�  �YS�<A|h҂�ѝs�P�� ;`�g[����2�t�����W��(ӯ)cmR��h�T,�Q�`,���N�ߏ �Y�A�M2Li���w-��|�����҈"7ư�9l7lW�)��q2��IFٓ ��
�r`�*y���;a�Qt�7Yɰ=���r��sl� kC�匓N�.g�E��j�v�&�74��3��Uű�G�
h5�?s��|-������v�+�,Y}����k�Ъ��!����.4-P�B�וC���n�����27�t��<Ժ��B�{�	�.9k�?e�y#�,�acζ�y+����Yh��z�\�yl��1���R�U���M̘�u��zN�ur$�~��G�!F��Er�yL�0͖u�y���	[Q�%8�x�+\���j�dBY��\��YD��I���.)#������,��%��87of�[�{z��|�ے��X�@�:M��	#�/��!�b/���Z\2��A�i���A���+m`�ή��;D
 L5������[cQ���ær���DI�vlUO���D���lP��R2u�fg?��@)`�pJ�8\8�\H�����w�VK{�&��@��E�A�m(�G���1M1����Bac������L��m$�vThX7V=zĞptOv��[�kB���(�b~�o�jk-\-aA\DiP�A��Iː�d¥傱VGeC��,rS@��a���h��k��.�M�g�)�횴?��1����Ž�2�l#k��q3k0�{e9��k\V�!�We��4��<ռw=����h>�~���-��m�B3*z�̟LҔ��� (�sF�Kk�N�	7���AU9#���1"�E�]#��x�${7�ҽ�Wz۷�k]E��R��4.	в�`!�q��š��43��:�qe@g6�~~�"K��&s�����4��e~�<F�k��by������pJ8�[�	Q�-ŃZ�=��i2�+2=P?�\T�R���\)��JC���s��|ݛ�%h� b�P����@2��Rk.]D�KYX�?�H��W��׸F���51���F��bm;:?n�=t�5^6�X�t�rZ� Q�~e-̚�#hWB��A�)��>iܣU=KVŘ+3�6����Ć^�h���Aw�y��g�T��V�q�Նd��]��|����W�Q�DUYF�����Ǌ�9���4�ݷ)���D��A���R.��ޖ�L�!�������/fܼ���,�aAK	q`HH~���ۥ*.xn|�&��_S��0!�,ı�9	���?ʤ7�dkk�X�{'�� ��Ą��Eov���g-���ʤW3��.�#gϖ\y��� .�,�ek�#W�$~^��2�d+�E��L�
��R7�h���Հ��F�Ns311DtN�ד�:�F�P"���rRE���*�C�v��,��:���ϫ�0h��̷1�
��pϮ���Ñ$+ԕޓ�s��#�Wr����A��6|"޲�iJm���
e�[���b3�N}�"�,�7�o��P��]�!��+�V���NE�CW��%��Ɯ���	��x�Ҁ�S�6+��u���:�&�"̳��� ����0��L��ri�_�io}�h��.\���ƘV�:H�1���R�f�qr�EJ��~��5�8d��X5�dO����ө	�����I��?�h���ŉ�D[]Jq{�K]q2�j������f�3�T�cZ=�~�>�^A��R�=<�$/``0p���9�#P�}.��ԛ�>V�}�7{�d�"-�-�k*�J����%/��������;�Q>B�.�zO����:�rs�ծ=������(�3�iJ9~z��>���ñ���;�$��Ү�B�x�w�.p&-���:0E ��`�9-m;�%S�hX�Ü
C$�O}f�{hh@��g��&J�w��a�ӆVJz�J�?0�ԛ�t����O
��O����3~�{!Z�@�xj'Q�B�{����j�����2F/N8x���)���(�c?�E{����M,��8����NSl��c7V�l��a�\j-�������{a�h�jC�D���~��z�����L�&�,x�}&hl��J���)+y��{�?����L���d���v69���7E42G�Ψ�,6�ۄo@Ryd=(C�V�E�.�r��&z�`En���h#8�E�S���<i�T�
�7I;d� �w��.��9	5㬮�:(ݦ�Pd�pJ�F"G�*�r��ʊ[w�+H�t'�-5��aD���N���iUv�?����J�7@�B�,]�DM�r2 �3�iQ����������.��Ͳ�����y�z�Bq�pEg��!|;ݯw�u�1�c�k(�X�||��M��#X�ہ��\P��Z�Vy&��9��6��X�}��X�rpZ��^��FG?����D�^rmķL��*����̆sw:��6I��u.�59�?9�w�50�eEF�w��T�R�q7}`p�U�Q�h����&[�(�?]pJ�H�MefH6�-̯ǩ;J��粮��Z��G�HS��36��C����gK+��Tez���h�LᓎTc��C'i�-�Y�י�D��A�!��:��1ń]�U֦.ۭq#ߑ�!�ˈ
ƥ{	lq�Ȅ��!�BYk����Ƴ�A7z�Q��qȣz�T��;r�Ɯi�]+'�=���J*W�/�KK�G*����DnBt��Y��R�43g���oj��_�����W�%�[�5�W������f�s֩�r��2w�J�t�=u�M�V������Iv��}i���iݢRj]lCm��ǁ���15�ܳN(@��ϲ	ȼ)N���ȴ�Ȫ��bh�����;��a�D3iK{�P�K�9N&^���g)�%,����q9����Iw�`�s�����٫p���P d�њFIU��si�З�:\�����|/�]��`��4�0�s�� j~S�P�~�u%s5c�uuB�C/c��nW���~*<���uE�m�Ѝd�' Iٴj��ߏ�B�k�m����8`nKq|i�D7v�$�/	:��sPNSh�A��i�fD��*�6~� �v�;���5�b��uj�`�k$�t���-;�0� r�5��Nl��3L4�G��!#S�ā@��������h!�[�q��x/y�Y�P�!ŗ]ʍ�<�8�j:	v���v�7����"�㽨1Y=)X��%�m�s��$�	�き��vVJ�[:��B�� .�[v��*�R�l Z�2����~C�g��ܿf<��v�#�+ݡ��^��y�*� �iiP�J"=7���ٕ�}�8d����ư�E.刮�|�=G�Rf�Ac;s�M4�� �q��<�ɔ0I������ҜH��>�֢Y
���ELFy��A��1��&٭{��^B���'�� �@G�(?0�RӼ���Y��2<R�њ�H�k���Z��� `W$Z�&�s~`?{'�o�>�?�?Q���B�4��y�Y0�)��%V���s������,��[z�^�"�?���#��^E��z�"3W�Si7Z�Z���t�X�T����C�#6��9��H_~�˿��z�v��H
j�J���bĄ��mH̅qa
��Lx��� k�Eo6z��ЫRTqv�J^sU}$�}-D�c�ׂ槌�2h�9zE�kl�$���WT��ıÛ"���DPo,t*���gM.��S����̹�@�9��t��n�@��8�w�������G�1��@��QN�d-jY��Z7�TeH���&��ˁ���ő��G�3���a6mc�^�Ŵ�MM!%S��>���[�j[��`�kzD+`I/���R���AeE06���21��D�V�mC�.�k���=������.�X�|W�]$sh��b�}-�\�`�.	L��i:�M�
�������摋&z�����@���q*�%�"����RK�B˻���AbW���-^~IeVI�$�iޏ>�o�m�5ð�p�5���kU*���C�5nx���^M�0�(he)͍! P�-�$�����?F�[z�tn󘹌*�M��կ�S�OX�O�  ���h�g�ve�u~I�y����O�g'%1y�`m��r�RC���?��|����
4� �Hs��ȫ�I\>Pv��n�`[u�&Bh�1!肠_ї�Xf/�wX�1C<�ѱӮh!/�`+@�z���N|�[�%��Lϻ������3Xk�@���[Nu�j��*H������+�j�>���2���Y4��"���޸3�����|N�-Z[�^hU[PQ���Zƭ���c��Z�U���Xp�r��&��EѤYvr:��V�[�T��:W�ku��c�^�y����`M^=8��j}v�V��/`F��XΣH�%�ˤ��>W �	8��j>8�>�B皬r' ��(��N�� l�� �|Z����@�v���_�<{c��k��#�� ��mO�1�z5vn�u$Y+'�h�h����� 7F)��U���65ed͸G�t��ou��su�l�pa��0xdx�RwO��/R\�YD�<��?��F>�1�C���:�}�P}:OleM��2�N�{1�0D���4�k?���>��2�z�,�W�yKa+O��=��ʡ,Qn.�3�`ٶ��\��4�UI�|��]�$����Ӣ�xFY��a���Xw�6��T�1���U��*��@��W�*�,�>�ٖ/!���O�t4�	y�ϴ�[<.4��kN��M�!���mI1�#�\J�qr���E)�ERPϺ;�<�V�����}[gL����Mڑ�e�ŕf�ߥ�gP�� �"��5g(v E���P�ϞJ7V�G�=�B�8�d��G����A������<��;A3��|��k�����O�H���g��D˃�����E?����
"Ψ�&�����Zi��-EcO-��9~���˱Z��Y�6n��ݏ�[1�۰#C� c�+�C�@{�O¨�:O���Im��1�mg7��v��j�Rw��1�-�D��=�Ttn�_�̓�P�鬚_�1O�>���D��ֹ��A�+���[��Dj|6޸=O��x��!��-�U|kñ_��Xu�Ӟظb�
P.�U��.�ѕن,W���r��g��"�A%y��d���'��3��א��(���ZR���e����2�gk����`����ʫ��«����.�UR�m�d����rl�=l��>(��iǑ�ƛ%���&)�_/�>�����Aʇ������e_Ü���+��N�p.��b�
�=�/�����4G0�C�&�Y��Ei-�P����Y�4q�C%��f ����s�_�}�dGc�����F�?1�,q��A9�v�ŷ��=?��_G�����^?<�äs�u�#bڊf�g��FA��v΃� ����?GY�@Zt�=ƛa,��@�|(g���Z3�>��m>�	۪R}m�?�rѭ{h�{�a<��`Fnڄ|��A^֊�E���QҺ���KN��u�`�dP�-?�_�z?r�# ي1\_ʹj�w��,��a�e��T��y�H M3bk��8l�����!�����z�寒�2�3����T`ͅE�h5�%5�$�-����m��yV���
��-
����
��6�ƩL���K$|i|d��_�m7��ʆ�E���: d�.�	��L$��\FKKc�B��%����MRm|���<�@��AY֛���B�|�zZ˨e��:��	�n��)��7�q���?5�,՞s���<<E��K6���%p���w�������6B��D��_1��y���P8�A��7	Z���^�t)��L,��Zhl��'����p��nr�f
�Y�2����Z�$�#����=�d!�Vr�~U�]�Z�����E`�����&�뒺�)�)'^�2�Ŝ����u
��	�aY���S�(%��)��F8p��ʇ��a�+�D��_i�F�4U�F�!��O(�,w�&�^��^p1C�ߌY}�x{�����4"T0]�@nL�ȃ-�Vd~�g���J���SC+h��r5a�<��D�	 ��uNl��(�[�pl���e��%������EG���r�ɶL�O����8G  0ѡ!�|mF�Zq|���Rƻv���D��}n��I#
a��\(�`���q�+��z�}�A�o�2�������rD�̺�7�Vk��xH�?t8����'���F������5�/8�"=�p`{#c���MցO��A'��|�	��oS�1s�'J�.�ґ�D�ƨ��T������&<��{D��jو���6����[�F�|��w�ꃮ���&cB Cw���\�z{���p�༆w���bs=�a	3/Xt�o�̘�c�]cG�����%����? ��������7�).mk�}v1=n={��8D�P�)_�:S�q]L��{J��
ҲKj5�L3�t�} v�87��(sո6U�z���x1�]֡���؊���ԝ��q�uV0	�<&��ǹ��#���Qz�^�G�m�\kj�mC4����0�{
��ʡ��λ�E�n�nI�3����S:�"�DN?n�|�2g]F� �Y�-V�&��c��{=�הn���pG����pfm觮+&�챁J`|X���&Y	DC��J��l��n#����<��Y$�+6Y�K=�-��ueMcoA�/qܭ7j�i��o��2<%���*�I��0f�:	Ƌ�Ҥ�-�R������P�7	�W{�F0�H��������UE�?Kܑ�$�`�9�k��z��>tR)��m9���iO$�ͥ�4��i��1�Q�ʀ�R�\+�L=Wߖ�*�o�l��m�ѡ��q�B�>O�����=�z$�xu�<�Xh���ɧ�s� �izs{.:xw��[�c4�ۡ�L.!uC	��D�E�nA����@���PU)ۚĹ��k�"*۾�.�6��w�h�Pe_�Z_p���?�=����
��/���sy|=U���&>�[o+ZB%�����'9f��s=�H�Nw�b�����{.���D�8�*�>��2�"Ҙwg_po��@�
�p�o_zXlxV64EB    fa00    23e0�����G,I��9�7���ky=��^�H�[/Q��<xjl���F�W���
Jث�DI�1�]&�Mapzȿ^&�e�����Ӑ���|?9ዅ~��1��2�a<r@�b�-ZL٤:�f� ��A=��fڌ�+2Ku�ݨn�~:ަ	J{�uvI[�ϦXӧ��x'��T`�W\��ٶ�Htu�  ��s����V��U��2<m�y��D�\�ԍ�zN������P#A���uł#�<$��#Tu�	�_��#��j��N؁�ɫ��u��T/x!�2Ӣ�E�5����z�����\͵u,^���������1@���WLP�!̏�}צּ�%-y���0�
9^��l2b�k}���!zJ"�*���6�(��<D)O!��������>����,H�N�J���	#�$�
��m�J�X��(�`��RI}�x��b���f@I�M=:9s��/�<G\��]\��Gtm$��7A�	�r�`�D.§�H��"��K+�'��!6����K�@.:������z����3/9�#�{�"=� b���(�1���ڝM85$��gS�軤K��ٷ}��~آ��� ��&��TP7����Qm>�O:gHb�e���j<w}.#�]�����=�M�'�\�	d���l��ZF�뉝�M��pJ��̟Ȑ��݃�:��13ʊ�\�*�B���ތ�k��f���-yÊ�u	sܡ��jBS$	�e��✒�
��F��*�]j.Z�;t��L�_!�iʅl�Ec�J��5�$���R����������_-���7L�%�.�}UI���I�A�vu���[{:�;Vr��V��%�	 �f$5r�V���l�1�zel����������䁳��v���'�m�����y�Nݶp�8֜N�ͫQD�HA����5����y\��Zo�]$!�'&A O�c���e}�����-�c������{~�4����P'j讙i��Fu��f'�ᨾ,u
��'ahM���vU���-�U��;<���N#2-%R�pL�Z��̯$/���6�P�7 z��JI�+�]����w��F��T��-V�{|@��C��wly���T� J�}��1��ڰi��y����[U/ʔ����qR{��z�Ȍ�W��yЦ���dW�@�![�G����jKt���RhvK��GQ-�8p*�����������nvK�'�$78��]�F��>�l^�rQ8�]_�r���(iu�xOo�Q?�xr�I	)����׫�p����1~fX�L�(��E	Jx�DN�UV1fAG��x��Z���d>,�}��D?�U2�P�C7KF��T�i,�s�̱��.�>6�g0|PC����v����Z�R��.�Q3��%\�(��{��I^<-��X�"���Y!�5��׳���$πE"���K���&�c������Z�P�c�S^�r����'^�q�c�[J�c�¢9�x<QِL�y�I��2���k�,�!�YX����9m���݃��< ��}��(�&(�y��Ĭl��k��#)�
J�`B�_��{��`�1lSP��:˜�D��)Z��ح�)�y��!�|)�ƹ�N|�2�^����È�D��`���"����t86�����e��CPG�Rz�J���U�.�V�A�P�eg��[h¢��H�t��(��%�A�+~Dߦf$�}�'�!��0��1%�N)IPm'Zl�"���R�b�us�ҫ�d @��9���Ӿ���q��HGP��#}�ֳ+������qʟ����Fl:�ɬ��rJM�'+�E� 7���ϑt��g;�J4U�X����M�橘2��s�P���7�d"]�W�����*T�'ݮX}g���}
���(M���n����&�N��h��U1����f(�]>�����'��s1��x�q�.o�������3�>e�z��q� �FB��X�Qs��-��9�s�T�����|��+Y���k���j�D�&�;d����h}�:�%['�O�3�5ꅊGț���Y�r�����]������ARr@{#1���`�f��ix�3i��տ>Mhe�hZx��WPlLZ;�Oۓi�Ϳx����{|"�9 >K�p�~H�#p�ː>��u�9zXЄޏ���w,ʾD��G�cP�H�h�`(��{1[���0B���M�B�t����@q�w�{�lQc����k�/�5�~I�О���k�6��Ն�U:�'ӥ�V�K3��&��<��A2�=p�$�f��p'���x�h���	���b?�xp'�?2 �,��[,��d�@@�+�3�f�R�~;\⸗\c� ���Uu��Ƹ��M�QE��K�o���o��t<���ޞn|�(GPt�����]IQ�z4R��gmns�V�@H��S@?�F���gK�q�C�(t́׹O\N(���U�|�]!;��:�O�sA���ޠ�̽ۙQ,pY6�n��<
�ڪL*�ޥ3F�S�>��S��k����Š�w�_�$%�tB{��o��t�^2A�O*�3����*Gc�7���B�6Go��W�g��n}M�0����T�" ޡC��xo��X`��:�
�ylT߳����*�GKxպݝ_��5�klp�my��׳,?�;KTf�P�i�G���2���L�Z���m��
�hPʰp��ҹmU�+���-��Zg������Bُer�
��#�s���[�� H3����{݆���rf��uhxL��C�{N���*���j������/^gQ��b:E��:�ՖD#��'͆���'eG� ���5ͿnP�L�ѝ��dᒤ��a+VX��oqA��޲O���W����P�ߒ�Xe�B�Q�V�~v�(�}_�1�����Y�B6��E�oX�Q�5w����]�SA;m`i$VH=ʶ/�e��n\ ��?�1S	}��7�&���������NC��d��#�~8�0�UN�}�9�#Ƀ�7���>���8�Ә�ץ� �FG��u�醮'?���1E�K�}B К�e��~���J%U���Um�Q]L�n��� �������z~���BI]yPE/nQ�}*��a�Uť>�l��#�DdL>1^��=)�$6�!�*�H�e?�Df	��>���W"6�\7vHf�e�����"�{�=��Pd p�|��FЃ)���bp����W��Qm%��e���ɟI]y�G4���fE��{ʕ+��V�i���biTINP-.��Ш��'���F	l�:�kl�S4ӿ�U�I�Xf
��o�8}X�K��X #�Yn�a����D�����M�C��),��e�"�,7�oZuzi��r��5Q-���8��-χ�O��ɔ�G;o���PT��5!��D�"(<!�2�"gwO�<�j�p��s��{!�m���y�q*?V�l����h�� U SV`-���ۣ%0�hKt&�Un� ��ɠS������K�i΂�m�s[�~=yK��SG�[ru����Ӳ�k��g�-b���%%���TL�5�մ�|Y"a�"�r*�]�.�:,��M��ޘ�G��~
LV @�l����:3~�FR�io��?���q[g��r�ԅ�ӷ���b�P�<����-Bl������E��h�Ǟ����[�������j��P����o���5�q#Љ�a�4`ʤd�t���j!q;^�0M���o}��
��eߓ?�/�ܝ�@�~m0�GL�<�SZG�$��I��H� �V�R��q%��g��G6�<�v�N�y߳ �sbC*J*Z�(|��,D�Ҽ��ĸ0�&hk�j��eU�pE����hi	W�'�SgZK�9��r�-�@��<N�����=�<ُx��r�����Ix�1��M�(���:�5Ćn��y�]�pQc{$��m��/��ԗ��=A 5�aLh�.�Y�����l`�����a����L�L9��:H���ۈm}/c�|1l���Y,����w?���;QXr���^{�Q'�[�=��r�m@�J���f�3�4�<�[b&�����ݠ����J	 �������]X�N���R��:�r$Z��ev��t/��5:9��OJc����J�����݂��x��H����H�DVTw�{�p|��șU�Kj��s���y���eTO^ϯe�NY�d�6��)��O�+W+b���|�fx�a�����NS��K,Hٹ�羀=(�OsW�x"2l��Ll��B'>0�&���+����Sz�$�b#.Gɳ*I"J\jjr�|��g�ȎX�J/�6���d�U�DU���9�Vk#y���N�5KF .�m%�w'�E��_Aؔ��R71��g��Os�mS]dګH��/0�[.�5=��hv��*A]�S+�fȋ�}�������]��m'���͹��V{T$��Ŵ��ʢT�ݥ�F��D�1w3�#|��J�_�<9v��Gu�S���}�X�S.�:V�6D9�o�����͓C�5&���mTiF�3R�J]�]bi
��S�=Ǒ*#��B^r���^�ySê�����#�z�H�G9ܬ|�M`�&��ks���tG��1���N�`T��9����R9r����a���~
(��;���f��V�[O�I�=�$�0���R�#2�
#efp���C�t��YwPȰO�G#7������d|U}˼2 &��9BO7Da2~ 6��M�Uޞ���jI�b[�6�[�&f��N-���2 ͠�y�a�CPm���+O�Ǥ�' Nl� b�
�D�~!�_s��x��s���Pw��z�
���D/��Bq�j\�0���G��&<Z�b��a�6���ND���ry�[]���}[|���+v5�&��>r���\?�L�ңD��tة��RtYQ͙�A��؆|j�[T6L�I����M��k�7�o��Y���YpC�.����_̓��8�'�`%i[nS�y�Xukk�����R��nV#S{�h����&S��`lӷh;�I�4����G�[VG?�yN`�f�Te��"%D�wS�0t����}�'�q�z,A�ؑ���"�[���?����qNx�����K.y5��K��2C�݆}&F����f� ��_ޓ-����l�\f&�2������L����}����pj�������rzo��4�p't�eg�-_��qL-�"߭$��x�y�Sj�S��dW�#u�p?2~�������"C�?���F��S:aS*�H_(Vj��$L܋�<�i�,J�V�Ukk���>�E�/v3�Rr�U *3
�Q"s <�s��g��(�{�"I����,7�)�рx��TyI�ľ��^(�S���]oZ�����OR��uJt@e�FT��>	m�S�E��{j�Cja�g��z�;֬/3Oꋫ�BZ��5���A�9@C�
9��m`�n����zQL�aG0[*Xp�ӄ8Я2SѼ�@x@13�3�\>���+m�Q��w5#�R͒O�e �S(���͌�fL�5bωȅqY����3�^�U��
3�Y��,"�=�4��&�7 v(& &侁ϝ|��iި�H$����T?����K�
l�L��>�-�����p���1l�p�/�7ɖ�Z΢{x�]�&=j��;�Ig�Wo��������(6��fs�������+4���2kg_�w���k��I�u��:��7���AP0P4���;��J""�^��i�Y*�{�L�G��:�?	J�u�YO2�z>�`l�Ud�JTjiJ���d��#"�:��|��(����0����M�Hah�]�ng�>�J�R4|������	�����<\e��jt��C�$��d�DN�W)q�Xo���$��n�8E�@��֌]lu�0I��;�b�
��_��߫�(ġ���8 	������0�#�rzte�
�W����E��E�������.�+���ll	�M��9 L���aO,;h��+�n�-*�m�
�N��co�²�����ސ��&���Y�Oi~b7>�&:*�>��;�jb!� g%���
o������_D���1-����o��߂=r,1@�+F�F�#��w0��}�Xj����1��ѐ/�f]�$#,�-�8��5H���?(�"xxq��x��N`ىו�<��<Osn���ڜC�&��w�Ia���EY8*���XS����a"FD��
��C?�ή���n#��gFp��j�
��|	�t�H�c��ISH�ucK>_�N�s%�53Mm��x�=I�?վ�x��G!UQ94����mf�"Z�j�'�����v!�W26�W`2UF���}��|4�/7]��A��̗X��(�~���E���at�Š�n�*��&�S��'�:u��ѹ��c��]`z=�;�[�%���H�O��и�:��t��	��ѸY�0V�A��"��V#"tH(�z%�õN�!����,�H�(a@�
9aEƁ �>	�fd�%�M_C��\�1JHI3hͽ�o�L��]ј�JH���%Q�c���ב�1bq�F�I7��3ݑ�.��M"�U� ��:J�p(��_?� ��5ImT����!	��Y���ݰv
������q���{����4��4���8󉸔	����p���R�I>;#��6s^��\��eiUv�>h��q����*%!�h�V/�H����'��6x�]��W�aX�/�VyqR��"�i��R�Sm�{�7$�]����p'5z�)��I�'0�?��Vh}N� =�ܾk]�ץ�+\d��<�YuM�2@����G��9���*���1�5Pƚ���7\Bu���R��?T�~�"�ïOf�S�!���r@	\����XY"�O�&�ф���l�GX��9�Ӗ~�������?�1 �L����J���	��P�|7�����dZ'f��Bo�X`sG�o ��"�=��*��.���.HS�gp�?-��������&t ���T�J��?��B�����kԴO���5��!��2ͷR���w$^D�/*ɿ'e�v��U���z�����)�EHaK%���A )�H����� ~dYЄ��UQ���5�S�����i����K��)�奛ѧfP���͚3�M��b����ׯc�� X@M��l憐�H��i�fL�]�*51�q����q���]���&]g��;Ć»�o���l�$���fj�E��~��V��Z@,|�qxT�߹ ��Nn4���vܘ3�Ap�X9n~�)�T퇾�>Ut�z�o��N�k_�a>KL�a�M&�"	I�فh
�*3q���Ma���1N_I��Ь�����D��T{�.��Ct1��m	��k��d̉��Rt�����79��\u�"���YӮ�}=���qK#F��[��6�#,�O��$$��KY&i)cK��m��쯨���3UPЃ"����r����q�1��x�y�%���W�݅Sʬ|�v���lDCUwU�LUr�c9/���D�5tkGZM�̐S4]%�@����������zu����Y��6?V�fzH8�O�M[S�a�����A�_��[�5\Γ5-�G=��r�6�+_���[�?vf|��q������u/>k>�q�/��D������K��k��x����K E�%�|���������IϦfFu8�e�b`_zv*�)yL�W真�}Y�_�<��
����R�c��=�	$��[�P��UwP�ėC��?�|�G9)�����h�8��&�����)tP�sg^���?z���5�zO�֏p�kn��OfQ_B���_)4�!�֥$��(���L �Ay'��������>h�);�M���q!}K"e@�:��6qn]E�b����c��ad�
���k{����q.g��O,umLmnܣ\R��][�X	���ɽ��l-����~��2����ME���tL⟭ǽ������]S%���41/r�+�K�E$��0پr�ݴ���T�\�Il�I�<��9���4&#܏i1x�sֆ^^�܍Qn����s9��^��a\�]�fB������M��x;:���5:-ӽ��#&��W� $��J's�A�Ӓ����o@�����F��T�_$���6�7'�E|��u�W<ypHwTV�.�(�ٔ�;�O��������`k}}�TIH���ĺħ2��+C�m�U�V�/`��R�-��"皋�q�t��Wzv\�Jd#�6���È�D�R#��;v���꘺U]Y���}�[z�^������=b��fG�oϼ]��Wx���|#��~�
eJq2��Q|6ض�����bHI/��ud�!�YZ�I�oVR�wO�Ȝ��ұ<@�ʀ��s��91�%��gb?`���]J0���N�U���\�`d��������~%�͊ڼ�ֽ}Ƭ~���)��B���eC�̏��B&б"�����|Q7[�E����g*Q	�Ƙ��pȪ����ū��ޮ�,4Ɔͬx�B�1�Q�wnu��;��aWLǠ�2�P}m333�6Y����_���-o��Qu�tw�fTt�q��*2��ߐҞu�S94�QÃ���}�R��N�a�XH��#��G�c��VS}��'L���cWf��N�޺�_��PY*��2bS��0Z�M��ҪU�T��`�뱌����m���u#����� @���U�:��AJ�Є��"���M	|�i:�`��q�[���L�L�gZ,���9q�o1�,�7"�P���>_K'�!ʹ��{�n��ٛbӾqFk��rRy�wZ��n�a�h��[�&1D��'���$�@�=
��W].G`��Ȉ�M�T���M J�%�~M���h���6N��aw,ߌ8^��K�Ai�ē�T� ��B����e�s�����1q=��Cd��GĿ��2��:~E�)>�he��٘���N�\	����d�Y{���I$��y߉4.�;�H-�?�V��S顇[�%��R��П�Z	�'�:1�lX��c�بS2�>e�&Ho�_�f�S:eV�7��"��26{&�XlxV64EB    fa00    28d0��
Lz��Z*��3�C��Ll,뫚i'r֫�~�)<w�8;�~+h�z~cga���6=�)!T_��3h�]��2��>���`yZ#��M�e�����|2LP�ZU��� .,3���R��G��+%���ѭpPI���L�;�ߵ�ݿF�ԌJ[,�*g}��&	$]�cź5K�]�	���%��(h������+� ]R�0������``�9���� Z~)l���K�y����M��j�+#����MR]�Kg^
��9���O�̢}Ŗ�%q�`]x��S�]7�=�{��TS���y�=�Qa���@��XN����'Ix�Ue�yC`��ko�\|��	��-VĒD�6i����n�m��ߐ��	����?rw�8�PF,7C�U^�7f�*v0W-2�����
Ơ��QVX*�^�~n3��%9eť�ՏfH)@�,L;�o���������#I����?6ϵgK�a��Zp��G�j�	�p0�v�����eB��r�ڹh;�nUZ{��"2��$�؜��%L�:�@�He�퐂+
a�&�Q���E�@Ax|�O$l�iW���a��hX ��)�b<��;:�,��A�_2����-���1q�j��o�4��:���j���9��d8J�k��ZM�F$�I_Ir:��9n���M��޹���@5E)$	�8Y��-�ٹ�1��>k1�iN'=E�}buY^�IM�������5~a�s�Qi�3B�p2�  y�k��7��Gl*��@��)��Y��(a�N�����r����M[��
GU66n�ɧ�� B��OM������ ���]b!�ݓps�yU�KH$�H�6�U��%��Lc�tz0����Dz�������H�^_��fj0�/�9?"�NO2��W�� �C;��!�DJ�fF�IgO"�x�dF��F�:��J�..'[F�bԲ���6Q������Jd��H���k`q*�i6(����p�Q_2r׵�*!�3ӄ&ـ�!�c�C7���D�b0�.��G#i=m6D1���g���s\KW�XE6��.���]F<�V�(����Tׁx�� ��ͪ�O=k DM��f.@�9���G~�AzT.�[4������/P:C t�����W'�p���S��h��,���ҋ�&1r���3F����$ͯ�"r��Vj��@o�FcR�#>�n"�����n$�d�Ń!v�x�.��ɓ�"pl�Xz��ڛ��PMN��^��ĵyE�!�*�&O�V���k��-/��@`���̧������C-�V� |��p������Cm�|ғ�İ^�!��AX��݊�N�OD'*W��`��TLJ�ߪ��
�ɗ��L|�����w`2��&:ԭ-)�W���X>_��ד 'ìc.N 6S�[� p
,_�IV$gP[�\��2̴0��o�T˂G��_��)/�9��м$> O�z�ߚ~?{���sC�(��KG�t�ܸͩ��.W�z��G���ޠ!>�i�ᙅ�Ҁ�$�ܮ��Z��&a��Y% t��9,�� c�C�E�젡�4��f�'��Vn�ne����t���J�S\\�E��L��V=_��w���j�:�>t!��ς���q��#�R�[my��f<WW$v-c�ޗu�S�U��=�u�Y@gq!-`��Zvf����-YH'�!x�m��f
"���n��`S���_��<�=���1nH������v�Ϫo�~$\@F�c���;_��9�ZśqxAEh��dg�s��"��8�Z��J�� �o[����/���i�yMm��bx˺����i�"�BN�54��{���PA��=Y	�*5�p9���C���/�������++R�^���#Q��c�{������T_N]zW|ɤ��N��dc��i��(9��+�"����"��GMA����3/�AA�Ok���崯&����^s!p�" ��Y���?`�=��S�X��\���H�S!�/1,-X�j`��#���(G�vaH�����4x7���T�`Ie1�x��oh���j�S�Д]�I4&
�G�yϵ2�>0Jq5퉈��B��U�Ϟ�:�V�6�V�@u���Ц<�&x��^�Y�?�|F�K�W��#��{FH�/�Abd�N��r�Z���&��
��W�j����mj�ao�M�<�⼯MMů}$�4¤`i�M���� ��|�Y��i��L��Bz'���G�Oq�B���B=n�����c���E�y/���c������:vV�Z��4�5P�D���%��w�[�8'�(��Zw���5�k�l�#
��f��p4�~5�����S/;�S����^rw�L����0��8ϐS��[��E��	re:�e8e�#�s?��S���[�:��Q7�z�0v> 0z
mĽ?U�۶�	Q��&��BM ����Ϝ��'�s �Su����(�>������D�A�-�A�ύ�HiV���Fj���k�c��3��ǒ�-#�C%=��E�'R;�ѷ3��j�e~t�H_�a��ۚ��jx-ҚV?J��"�͕x�U�BR��MڟN�% ��'ك�X�>�N6��H_�a�n���ޭs�6� �e��!d�K�[،�j�f�x�MF{���-���Pu�
8o���9.�$y�$�G:�G�"Z��{���3v�ȶ6��>@C(��@hKt;��v6��Wtͫ�^��e[)*������1͒}�(������g	(kþ�9��v����:�u	�q���?%!s-�'���l&�Ri����0��+��	�>���C��reҏ�R+w���T�Q�k�]7�m$TEs�yJN�~���q���P�RYV,�0�C��?��͆.�@������.,z�t�V�'��sW�ӕ��Ɯ ؊�����ac��a̿e1�|1���6���u�b�L���)�t_��
�AL#�&�����G. ��ds7�96X���+Kr��B�Z�Qɮ��[�E[��U�͐�ő�@�DꖜF;K�Ķ��l�=��;��>�?�P������e�V��I�6�����<�*��N��Wɯ�q�EA��V:�[JwK~�"��q��D��d�'0�٬#��7�`*���X�
7)����.�y4ץ�]:�;����w�s}�߮�x�ޥ�ٕ��Bd�
�n]�$O~a������*P��2��i�o-H��N����	����'�u9&�h��̭��O��˜<u8wH������Z�GKt�����i�γ�_�8gK	��?f�:Rགྷ7��Oh��H)�;0l��W�u��'K�tjqa�oIY�n�Ľt��e��o�>�.���t<�@�Z*���[�tP�������Z�Y�d)򵼷��p�����<�/�KItn����Sh�����%���p/��c��d���x�p�g5��_7XZ� ���)Q��6Ki��������)��r[��}c:^��U��2��������A�J�5�g��B�Z�Ks=�d�p��A��6O8��ʓξ��7���Z.��W����=k-��q��,�� x�w��������ceX3�y	�H��׬�rx��E�����ˆUB�Ͼ��?����"���ʔ��}6�S)�������T�x�r[�\�!�8u�#]+b�z]�<��?��Y;�N���J�^��\f��m�@���ƟRp|�ע�3��O�4�D6Y��S�˭���)D�/�a���3ʖ,J�?�H���1v���[˳3�s iڥ[����x�ixeK.>HI����L�H۸�F���	���3B�/���'�V�˹߼�8�D~�����Aq3��үH����kOVFu7�I��Zm����o̼�V<�`�e���R�A}�Q�#�T�-M§.�5�?�@�_ƪ�<>�h1���F��F��uX|c$F�S��MK���Y��Q�`���4���tOj5EtG^����C���G}��ݛg�˫��X#����՗Z GE�OL;2��ۭ&��D6[�J����I�F����&��U>�8�����t�;-����.R������#���\��� 8ׅi�D�]炤x��w94K�e?)��;��;�F&g,��*��MY�@N�0�j�]~Y��ƥչ�B[6f-w��צ����P$��NP��:J�"��w0~��inxY�aj��8�T~��g��������/�.13�����l_��J��`�)���*��C�5+g"��@�q���4 �W�Q<H4����~��戞Ǭ�j���jC��3ns-�`�.����c��@��S0�ܢ`(.�~���+��H�[VE��'Ҭ�.7��(1_�im+��&�ԟC h�'c4 D���*^LP6��w��SR��Z�Ѷ,	�@�qS� ط��?w�{��$n�Uk�����:޹?��[BJAQ� z��^�j����ۡ��q�� ղJ�#d�E)ska�l��lPHQ��m)Q���9�P�Ѷ�.gZ�DuB�O�����§��fQ�}	Q���j��8�(/\�l��bQH��R��41]�U3&(?dD䳟�g����ʒw��a���]=����M�C5lM�T�����e�<���R8ڮ/W�+�
l%�T��Q���ʔ �@N���s�O� �/���4X��z؂+y.�`P�?
��u���u�]�:~�����7~���9��l;=ܕM���;�W-I̐*	���{�Q�M�)< Z�/ƴ�YoZa�x0�qg�k[H5r��fR�k��fb"�y���oe��%�$�v+H��o���h��f��;9�@>̠ �~�g�u�N(�v*5��pކή�فZᴈ���؛��;:�g���]]u�:���*j��C�{�Я���G�w	a�*�
�����{��P`DM�6j�����5���jd:w<G_}.�U�s��_ �x�0Z�)���{�]
?S���l�P�����厸��"<�5V¡Y� I�f�J��H"6�3܇v�M��ͽ�ytΥ��Y��&#��4_�z���ug�#�E��Y9��b��E=ލ���7	0MhqC�̮γ�P�0<�"�������H�"u������͟����p�	Ϡ�w���i >�ͼiא��{gj�0Y��B�Q!�]ȎB� -�{���۟Hkf|YmSY8^�1(;�5�(��x��\;e/����#Zh4{�>0�)Zk4R�#x�@!|���鏓��/Y�N)-(p� ���|�q�P�vȺ��4�	��5v�<��т���܊���3�qO��R7�V��Xp�^
u���p�:5�͈;����e�)'�$ʹ-Ok9{��W����%4u�4LՋ咮鰿���W�A}�6fj~W�v����E�V2�ˈ`���/z[��Mrb�Mu�L9dۗ�.���~T;ls�be	����S�8}��6���J����m��֔<j_\أ�\*���Ў���!f7Z'� 5���÷�5mCNr[>LUX�N�!���V�m��݃��9k����6��c<��\���"1���h���N��sJ�J:+t ���a˱X��`���w�!�Y!���*�$��F��F��LF���]��Y�.�Yk�N�0q�Ȓ�O(��#�(e��qrŁ��8V����I���3�^�ѹ�D(�_
a����w�.D��4v9�k�HD��q��Yp�-���Z����7���"�m�j��1�VT&��q�,)O~,C�U���/<�!3v�o�5 5<��
�)��yR�-l���W��}�x���ڬ������H[\��
�́�G�sQ�/�CY�3�� 4��nHX2���y\u0�* ��Ef���
���2��DRW�Շ#���U����Ց�W��6�
�%�8��L��XjSnpN6���kmGv2
�j%�v�5��I�L� ����-�9-y^t�	�I238�2I�k��>�y=��Kj���h>�;:�A��`�U�?B�&���V��˗�1�e�A���� ������S+�7�"���`�PF�uz���g3盕�&@]+ӊ%�\gg����Y�0՛��"Z��������Τ�CMR���怎�%���G�]~�1�b]0���}�tJe�t����U?	54� U1���x�L�ǚC!O	x��h�gb��J�[:�6�X\��������Љ��LbEK��iј'���T�T�<�	7VM����R{c��Z�_�,`~B"����&��S��\J0-9y��_�a 	V�Xk3�$ø��v>H�e��;PaS�9 �⫷9k���^���ߢ�?+b�^v�Ҵ��b��
j"j$�v\��q���a�`��%����h�^%W���D�-��%�«Y�5qB,�T7�ul1e͢gN�	1���s{����Bx���ۄS�,�3=+Z��H�(���+Y������D�E�����%��P�������eƧFSv�� �B�W�0�B;U�,����p������~	��S� �ӻz%[IƼ�m���Vu���۪L��4;�5|L'j��^�U�$��f�����6]gv��T	��<��W���7�	M�Z^�d�½�1<Kdr���D��dV�D����M����0��3ܰ�\凥-���/R��PFff��yHk�d:�%�4Y�0�O�ܮ�E�u�-�ƨR��Rvޚ����|J���?r#lr����q-��t`�L|�K2i�J����@99hL�Ŕ����v�o�`fo|{A�*PzG:ʆ������%�w�K��N�5.�{�rh�s�-�y�A�L0��2BH�'ւ-bݵ���_��z���Ұ�g����kH OFr��7���v��������%�:ѯ����IN5��v�,[o�ִ͐48C[�)�9)j���C����ˏ��	�x�6��=R�YjpCrŋ��k�*;�y��S0SG�6h�Rb)�oҁ��ԦFTH�Y��#I:A�I� Φ�LM��R>},GZ�o�#�@�4�X���8��_W��r������m['3 �6#�h��G�:Gڳ��F�>w@��YFA��T%���Sx|/����<R���ɦ�ŧ[���@�K���9&/Z����cM��ղ�~���D�������ìQ)��	�Tb�S5{���ƻ,���T�6
ctN$��	�r�ZA��(��<����%��E��tCz����$�d*-��C�~!���r|��6���I"�`s@�c��:�Ws��`�L2K!Җ���!ѩ�� ����1uZ"Ez
(�H��!��{c��`��_����&��U>t\9�ɢqC=1���U>�q��9��{ &î��L8O�D?Se�Mx��_�2��<��J��i�+�)�-V�� �x������>�2���sY*�&�粲C��2�zrBb4�i�T`ug�M�+x����9�4�*ی(�;��nk��tl/����|tPV�H��08"�D)��:��Y/�n��4js�R~�a�<�����2����'��$^�aw»랚�2og��S-�&D����FL�{�i�����6�t?4���?0?��1)���UU�Y��7W�_P0�f��Y��`�1WU���f�PG!&v�}mz�k
�/yl�N+&e�m�Д��h
� �{��ډ�0�4��H\o�5K5��P��+j�%w�5�3�����Yhq�R��o�����?��f�bѧ��r�y0����M�; �R�n�����dU���e�B}��YvCD�� �Ӏ�Q�:K�_�!�����!�Tj(��a�S`w��i�,s&��p�"���4���!
	-��g�7��v�,�hp�Łq ��s^}�G���5;�TU?('1'�{�����!;hH��
�G�I"+���"0!�S����I�J���U��hzi�]�a,���ˢ��U�lO��$���7&��i�ox�%i
�b���X���s�Ys.�{2G�S	�4�J�.#f��"��x5���G�h�,�1�M���p�;�F���`$%
E�YDOX�ۄ���$��D�s� ����\J\]����4���6|�[��Lm���2:�Z�[�ɶrPKGN����kV)f�ZI�=#k�Y�)_
�/Sg�L���MgZ��Ǽ1Y �i��ϵ3gؘN��{쏎�fP�����t�Z�u�9MԮ3�i;�L>9f���5��Y�Jk{k	�l�|��[!C��$�\%�'K�Q_�6���~,HL�����ft�`�j}���u�*�ƚ	v<��{�v�Y��0!o�lT�c�ZV�yx<؛|����`N"ڛI�n�s�ۘ]4�]��0CZt�-ʠ\Sen���X	)�K	b�s��3�t�G��Pp;�����|�l�L�5 ����@y^��U��ˈfV�$�~/hB�U��yIO�e>M�2޷v(��M�}����b��HC%�k��ic��[�<Ƈ�E#�Puk������т�ψ����}H	l�Y�{��#�<�p(���ļ��lA�+���
�c��֮�[ϋh�������ejf�#��k	��<��"�t5.��E�0|΄�4�9������S�[AKv��� �>�����SX���sߨw��_ wq���mKO}﷪�� -��ɷ���*�o.�ʧ��䤷����b�`��zw��D� ��-9��Cj�i0��|�\L�����|J��a�C�(ױ��䓍~w�r2�*�����#�NT�fg7,��
����EO��M�۔`��[q�σ|���t�3����]��\k
7�E`��l��ie[$w:;8KxL*ޯ�9���o=��L���mK�ak�,�<��^�R	�Y�Ut�FP������%ԣԎ��
HS>3H�*X�|����7~�y�I4��'u�S��+�Iz]��!���2CP�r?��EgߵJ@�F�_�d���y��?X�A����Zv���rI�-$68�3�
JR7�JD�- ���:���$~�����7g���j���4A��%�giHR��8dv5�T��6�9��6y��tw̚�[MG�A��p��6�*���W��!�s�#���޸M�)�}�t"KPs��e�w�ݢaw�\Ҡ ��Y�i|LA�S�won�u��H�Ϛ҉"�c�]���w��"����`��oO8�̼v��1z8(��t����}��7�/,R��� �[y6%����k���G���6��c�qJ�|}v4�Z�{��4�����N�VF�ua�~�0!DG!Z2l*�;�p} y�צ��-8��X�u��š����'�0pѵ+�0�`�X�HH[i���~�H*/�M��'���q�X����-���f��^�:�j5k�4mڧ�P���B�/bb�ƌP���A@���󩑔� �n�&��S��\����>�'��m��.WW����_�>�4�q�Ƙ��p���VV��]%�ј]�M�h�"�>cD ׾5�q��ɠ����a�4�|n�!Wn�a����W��Զ�m֧����mrἶ	btΎ ��'��5�T/�B�����'|(�Z^��iDrk}���?K�g�c	�(ɰ,֞`�)5b��	��_W�8�:֚�Q Š�2�E���=�r�I��<{��D ޒ?y	$hΝ�8���)d���Y�j�e8vX�i�H�ĖZ�7��!��}��x�?p��I����vMBS�P1Ϊ�=et_�ٜ�f�\&5I|�*1|ˊ9�`+���PU�iɱȁ4۠	��=T^z�����3Qʾ댥
���lt��c�I�&o��+V�8��7�-��3�G���u�qm�'_���j��W;�<�1^Ej��P ��"�9�H��2׀��?����]�N������� ���g���4�i�ix��q">g|�Z�%o"���E�y�lV�ۃ<𩺪�Jo�	S�k]p�V|������S����&4�Ѭ�w�?�` #�E� B��"�"�z4&�8�,��\��N�sî���o�Dޡ���S�D��Q܌?�P�����k���N���lp�l�k��T�w�iŚ0��Z�R6�",�[��?�{���R2����+A���_�Cn=��O�~���}���+���`���Ȕ[!n��3�P�Ȭ�eX����u�+�- ۢ'�6��'��%�&\��{RSѸe'6�EM�������z(����|�NS9�� 9Uԝ,Ͽ�c��g�E���ʴ�tq�n2S�>=)��dD8�W�U��xߘ��B[V���mcyNc���� �v�(�����?��_X�XlxV64EB    fa00    2540�y$��O��%�t��w�rd[x:��ň?�g���'��XobFЂ�����h��(HG���5���4���ܡm�g�dT;L�j�u�t��J�F�L�*�w��W4��+<C�&�����7��^�?�ѱ��6ԸH�tF��ܳDf�3�=g���A�)��ݔ\�*$��!y�/�c�R�e`��,���q��FjEm��{���q�xݿ`
�}1J�?Ů�5�_�(�ý]@�.EU���=q"��<
(�-w��%���	<7���z{��?�l ��1qň���o2Hcv|.Z�
~��E̝�m�\r������9�Rc��H�3�kм���*r��]]u��x�<>�kr@�/Sè]��]����|��N���+�xl��.�w����-�ķQy�ߞ|>��!B�^N���ޜ��f������R!�|F�8��>����ˌCq�*�!�0����R�LB�ElJ��s�B9ޞ/ӹ�P�:L�
�.�ߣ��4�6]b���T`$����yh��X��6� ���>&�g�!��R~�!����5�ӧ��D���wN�̛hC���5b|��%�n.�"���7�vUYj�� �ud�G�+����qpэV��0�1Z0.ڮW0�>���
�W�۸Qn��[�G,_�3�����F�4�Mp�D|���eh�)�i��?�+�m��TQ	f��-Y��A�	�B��۝O��0��<�|d(����<YG|@-���us����Lk�9�+���@qFW�^*��!�)7�3֠J���4��G�>��Mm�<�y�R!g⛉��;���X"�s��I������܏*Q���he$����,V��^͊����a�"a���!@C�1�T�1y�C�rV�E�CY}ٜ��W  ��>H%��aQ��৵��nl�NK��,?���CJ{�D�c�QPs�v�Ɩ�	]�a��n�Sջ��;^?���Љ>�3�k\u��wv.ٮ�Ҫ^�ۭ��؄qj̺���[-K���䪉u�`N�*R<��wo��3?n{gL���s���`4!<�*M�W��R��"�3e4X	O�D�X)p�>���WD!�07ʭ`�L�*8#teۓ����p�`�hq�U~�E&]'�N�t�w����q�
N�Z���
xR�s]a:nsdk=;a� �^=m�.�x���麗3�L���Z���f�o�T֛�8��g����p���9]/Q�0��F��9��x���Eٛ �K��͑���	s���443�`��"�S-��PN_�+�E� ����X>�k_��c�a�����~��7���v�����`����6�$�{c�o�b��H\l�5b�Q�/��o�����vDW�:�|;��������J�fM����e`	mHу$M,�W*w�d��9(-=���
�d-$�� u���L�8�g-h=N<�b�Y�X�ND��P��m&I5}��{�7�._"�"�a���JTF0�N^�ZZ��Kgh�8~�8�u�R��Y(@�f�|2�����������K�FF��:���'�- �a���v�U-F�H�Q�[S{�H	�='�}��.ъ ٠� ��I�?���΋�*߆�ְ�%#�^U��,m{��+T���nޙS�^g�C�i��it���b_%J_8�M� ��HCm�k�W���0@�m����i�N�QV)�� ��d0���r���{��2�k�89�����ʧ̓-���nC{dh8���W_��Fj�'���M��׽��i�����n1u���ܼ�+)��KAQ�߁|�˅�t�h/6�ajڢ�$�I�KlPqțb�fK8�U��f���2�� ���S������[Ѵ[g�r�G)E�ބ���gr��D��^�_r���5/U����,�v̢β9�.������ʱ��~�9|y{ǜN���_��P\�G?��;�����Ssa��ߡ��	}�Bb_�ѩ���L�����d���w y��ۭ|l��ئ�e�v��%��F�'icF8�$ꥎ�az���R�vӉ��o�ZD�|F����	�n�c�������ʃ��G!��}C�{�6��fmq�t��߉?i.%or�7�[.�}S����[�+�)�lA8;YB�.�Z���+r�����v�D1�5'���c�����hy*��el7-F�G�/$��b�ӆ"'?�CX�%���fs{&8��eO���u&&5Lu�.i���n���9���ۉu��g��+K%��aN��x�����9��gI�5�&�^����y�1�C�9S>{=��z����8@�wH��(e�~p�ꏋ��4�fɜ4�X=d`Q�(�O����e���6���Cg~8��������a�g?��� #J0�)�a�P 
Ǹ�M-w=�^H�_ڪ*�x^��P�~zkU7�('�RG5c?�r���
Z�v�vK��t>�]���S#]����}���`���ۉ�:� ��t�[�ӤȲ�f�g+*T��SsդRH�SL�l�I���y�wH�e\ؒ`�ؚE��d7u�@X���3����#�/��;�P�#&��H��D�׹-D1xo~��fذ����I���I"
����`E���kNd(��@�
�����\L���1�Fl��uÌ���!��&!V��ZB��Q@R�{�,��^#�m�, L�ʊ�P���=0��iA�3�}]����l�'��:p��:�c��O]�]�X���=��<|�X��?`�}�$��ː�	�Ts��L��m��(�5�+�-�^��p���~�eH� ��PBn+�^��XΡ*sYL�h�Ў7���W�*��l�Ok��9Cp-�dmۀ��q�wjʎL���α�O `�O>�Fl�����{ H#;J��뙟��e���}>8�ywC(H(��c�]l���w�'������5���=��e=��4�fݼ��Ӥ�����ڧ%�6��5�-��ԐXH��"��i�4_#�\Č���.ȣ�h��N_�2�"1�W�=[�*��p�p��怼�������� 1��ZI�O���s�Xߤ,C�c��4��w��s�viR���"6AF`�
saB��fKl�7ʻ�)0��ç��@��tO���#>W8ty�@^P7v#x�3N�.���Jo��G1��f@�����v�0��+�eK#Ț���n�Q�[t���Eֹ}!����{�8�X$ň�~��j�W�Ԅ�W&����S�7�?kϢ����cԗ���O�K��,�n�nZ���@}$�ؒ �4`AV��;�?��V�X�%�maLǮ��yeq3ؙ`i��<o�Z�馈�4[��Wr�z[�����Z_�Ȋ��g�)���ݪ�q.}���*|X
v���F�/'���Vm�{E�֝�F��M�cb��2��� 0(������"-�:�,��r.�r9��D��g��m� lBzT�Ӯ�e����!��*���`=D.����i%@-y*�/��7#�C�!awx�����Ԁ�\L���ܹ��w��E)MQ�a�Ug�U��
�_�z�o�"2��"�a��jXWHo�'W�O�9�-�I��.7���<��U"{����%)XjQ�G��X��d˂���S�Bj�O��:S<˞�J��ʿl-��y��� 0��ȕ�nы���q��Ug:�mw�73�=�Y.�@hp)�x� -��+S�Ęٞ�<u��)R��B<XJ�	�,?CF�����i����E�B�q�HaV<vX�WԾ�R��L��4�|�|d��ME���9��uWݹ��/VӖG��u�I�'�(�n׶���/��]��NX�<#y��//:��@oS�\�����"�_(V�
���v�YPhL l��,�Ծ��e�o�x��2��k9w8�7,�6�3'Ȓ�����V��Q4V?�Y��XQԛ�]�(����:��U�x2������E�Ȋr�˅I����dOi�b[���|��M����u�?)֢j'��qUG|��2=��&��Q�E��'A|����֟Cֵ����p�����ZS�N��<ev��F.�������b����=��x��D:��%�y^�D�C�L"����k�.N��>�����0��JV�/T�R���,y��W��ީ����
�~�q�b_�W�h"���Z>�����B@���LS3(l��������f���S�������	�O����B9��2����hFl�1�Ś�\�ǡ�ۚ�XW�~�r4�+�Yx(����/�tA}��0u�>1�O�;[;(R-o�gC@72yC����n��7�N��UB���T�@Fm�hnıY�������W������H�"��*g�!)��l���9v�v��zD�ΐ?_�-�Cxx��T�!���#Ս��*q�@�5*߸�d�� 𢺛l{&{.)��<d�zi��<r���"2�.�w��t�e������% ���I5&�)�w0�X<�ͨ�*r���ӕ�����!��>��*V"����z��� �({MpԀ�*`�X_��hw��&��P�~o�%|VfKP_F�-Di��E���(�2uǐ���<r�s�����f���w���y�44�+ؾ� ש�-��0���i����,Ff��y���GH���wI܌x��`P���Q�'
h1y�U|FbP�'!O�`Ĭ-��Q(�m\+���:9|�#es�pᛉt��z�ŭ�"�soyڶ�����/���7k�7KS)h.ԟ[��%�ϱ�"Ƈ��>�G������;���15�Ƶ')���K����^%�AB�f4h$ �mj_`l;l^h���˻/g��'�㦚�0��Uj�ʿ�+��IR� ��Ӷ��ݻ�8�#�
;�'����@�����5w�� k �LE	���}S_<�[��V���e4�����&�.+�Q���~4���RǊ,y?�I1:������+�r�;���DbO��K�[vno^����Z�2�z��z͚hT|e�:�)�v�}��of��R?	�����懾be����]��&���)tW��*S'y��������Zf��)��ޑ���͚���a$?c���b�E;z�����a`t��N�4��y�*LVs����������cH�p�]�|5�mƿY���^��8�K�x��JK�8˛`&�d�`���Dϔ� �����xP����kX�E�����4p���iڃFm��bB9ӻ8c��co߰w�+�'y��͙��;f���!�!
���`����J�M��{����"P������&^�;�����!�:�2S���&tJY�����OZ��$�W�8l�[��5��t�7��,]�_iJ/�����5;K�0RŊl���S7��?�ʼ3��{�7�h���O� ��OCپPȘ�Wl�Pb�	\G��4����[�7$�+1h�0\!h~����KH�2Q�3��A�>0ʚ�ʓU��N_O �n���O�8�	��d�/� �� �=�����\�Nar�Sr�0h�D�\"<�`��쇡�
maD��e��PQ��������Y���y���gZ�r�К�e�@� X�bu�I':)�k�'6̾=.x\�(�R�''��#:˰xy�^͊,�.k^�_��`�?؎j��3(C�h�;YpA�Ɔ�.2?��O+����œ��kK��]���Y��ga�t�x]{U]e*9�?[U8D�\�$�;��� �L�7��(r�(��rL��n�l���J�~����-[��{��Y7�<�\**����Lo�_�.��A5���Ƴx��`#B���@a��GGڅEe<�Q���Q�-�CB@�s�4��Z��k=虣�ٛ������5$0S�|,��?x<�%*��1�=��%�Ѵ����L�_�\�D�?9��䏆'gĤ@q���ihi�S���@=�F �Z�����Ȁ���k���Xj����ܨe��4=]��7��a�A���\|�[�����,�z�X�?�Q�Ƽ�^d�����#�z��Tfx/�B�s��4�@vX�.���m>��L@����A�����5�\ᠭ30�ڶ��g(}�����B���~��\���8��>p�a�2���%-�(`^��G��­�7y�$2��{!f����m��W(�� �*$jl�?�&}J"�˩ �m�"��xm)̐����'����o�$T����>�bT~}ȱ�^LObh���e2y�(R��Z�� X��+����B�}B ����r�\y|���8K(�����$[.'h�t�RУ���A��BLx]o%+�O@�Y��O-��B���:���C�5��C������W�"�<^����g��С�yAAP�m�@�Hc���DLZ!���`���Ah�O�Բ ����!7��@c�j�!޲
a���*!�,ҙGָX35]�K��2��������x�U׃���;��稏4��#�+z��'����303�8���}�X�x�	N��iQUiO(@��:�L��Ok\DN��\d�7L!4�s�K�Wu]�Af��tLYki2�-Z�5��N֍�~GnN�X�����*��~z�k���8�~�b[�B��4����ȭ~��
����)<?KW�F/�mf��,u�5�i�Ta_Lѵ�F�",EC���5��s�"R�[����C�<�u��%��TI���U�=0�7;0
�O�?��)�T�ſ���;Z0���g��V�������˟B��AɋO��5��	3@:,s��+�z=�^R'P���f��vma�ˬ��Y�帱�2h�SU�����ܫ��Yl�V�s���!�;�!W/���##�k��N0�q�Z�nEPi���/J6̱�N������T>u��������y;�r����/�=K�~(���m?���i�ѥU��ꢰ"���=G@W�u
-@~�b������N�ޕw�ײ�&� ˭;o��](�6��~5� �E���99?�?�k3��z���|�@�e/hD�
X4�I:�ˉ��Vf#;���l2�x�!f
�=o_Yj�⦭��
�N��e��7��6�������'�k����B�uA)����6`��Џ~�w����?��=I�y ����#oT�~%� ���F/C�,.�;��L�5�ږA�;��)ϳ�6�Q���e��x�^/�>�?�8��������{���ǰ���O�ɜj<?w2͐�z�Ѐ�ݮe�zi }X�P���f2M�-4�
��qۚ��WJh�qe܉�;����j%��E��c{��|�G-?��Z�?g�s9�)� ���H����(~�'��=�W㪳G��L��O6��&,�sO��@u�I,��K�^���o�����'޾[��Y!�7#k��o�����,��ᙃ�}��u!4 ^�r�@;[��3HP���%���0h;m�f�6}�+�$�g����8�@���������e���QC�6Ē��HZmJ�1���њ6<!Ȣ�d���/U�6�:�})v�=��֧Z9�L�t���O3ݣ����a��\�n2M�o�cD������� ���""Qi��ۆ������J�Br�x��!�6��W�dG����]�:��5�&��廛Kɱ�p�s\�3����$��`�����d�A�f6k �D��l�]-��l�l,�R$�gX.L���Q�(�s�5�`��,�/�.���m ���2��h��>
.�0��E���H�9��6��������ȸCR��%EP��z���1LwZU�mTp�Ky2$z����RWb���Q��NU��S��F�^}j;i��z�J�����܆���g]u�?k�UK��g��ua�p�
AbQ�w��
z%S�^ޏ�#���v�䦯��|��>&����f�44���&`�+#:����Y��$�/u>��S�����I-�������9�*�|U��&g4��(�&���Q�/���z	C����#���gn���A�F{������N��F�/�~����7]��A��q����U#ʸ�U�?�v������Q�韔��
	��u�5����׷OZ�^�|s�&��=u�=�:_Dm���輳߂b i b�1o&�l�Hs��C:�~��y��E����~�G|4Hث�yR�!2h���x�C�
��7�.,���Vfԙ�����K6���y��蒜P�T -U4�Q�J鵤���p0ӝ�07�e�y���s6N';3�Ɛ�?w���ќ�n��'J,h	*}�s�݁�X�z��8!|G-�p��-�� ��2n�.n�ًbIv�c�P�|,��M�	�I�G�sm�APeG��a����[��ćT�:�\AmwH| �>H��e����4h�y�*]�-��l��P���+��%�`��\�Q!���b��T���m>�6�"z��NdU9�<�U��G2J�}&��㵐4�Ջ.R25O��Oo+����`J������`�|�P3˄N�c��/L0"���j�bd�%�ZA�e�箏�2r���{�-��c��+&롎�����I�8+]�.��\I��m~�f���tQ\0�*�1��'�B����)��4}:�쪧[ywa#���hO�γ>�����
�Em��5�͠-ͤ�]���]ψ�׉���hU/����Q3�#E�	�R��<"bM�Auܚ��������s��N��� A��S�ɢnȎ�P�Y!<��v��(o����H�wG���x�r�ҏW 6|�|l�Ys��*miD���R��6�teq$p�I&������K�!^k�xj��*�R3�Lv��eu^4}z� �S���ɵ��q�e0�/�	��)��F�{Rp��2ݪ#�:��W�����wW_4��}��UPf����;uNOn���=O��Qb�����h�P��ÙC5`��l�W�"j�Z8�s��S
��^���i�h]�&��q	xuF-5{X	���դ�iS;��:7n��G��i�h;2�.�wU�;�s��`Y^PQ	2�*1 ��;r2Ai@_"'�8���ܒ�����F�&��@?�oе���|�%^��Ey���i��H��e����aQ�k:s	�*J�S��7B�<ɼ���7�m�a�iDd��4����B5�e��#�۟h�g��_Cqp?���A�KM�:�V�<��Z!J���B��r	r��Y(�P=bݵ��㓮A�EE2��D����S��}�:F������!�,{���ח!�aDQ(i(AB@�b�R��E�^���T������~�s`W��Ə�=��n�۶\�lӨ,��<!�� ����Jqm�5Q�F�Y�'�OL%!��!�\A�<{$���1��qx�$@]�D �w+�[Z���g�v��5m�v*Mv���:�`�"F${R�f)}�(�Z�]��-�B!0�k7��ݱ�����jkks����XlxV64EB    fa00    2600��ȅ�p���G������y<i�Gt�2nf.�	X�O儒�}�W�a����Kok��;-��ma�V�'�֢p2�"&��5]CF���T�[����9R��:KZ'k,Rb�9,@VC�}�v1���}7���Gu��ގ(@����8ܪ�S;�ǩȉ��Ȥ��r��������ML+!��L�?=.�v�aY�e�;���z>�L��<uؒ�&��ϕ����;���r*����Z����k���K���9�cj(��/O:��U���wM�ɌS�H�	0�Ƌ�ӛ�|}��k-\��{�c;J�@�����c<C��- �Ȗ;g;�@k�۝'n7�#sb/x���"O	��S9!���\�h
���9.�R�r$��oF�����	�W��͸���N3!��
��PrE� ����n-�ۀ��NA��_Dj�R�_\Sm��=	�r�c�y�N��\iQ�(�C��m%����|=܀
�b�m�ZS��p���
w��ʆ�O�!�#��jGҡ�c	_sa��Ϻ20�syT;��[.�h�&�ʯ5�9V�1��a�;L�"���,�Ll�,>�1�G�am�-�5`x�^����O"U�|���߿X�i�)�=�C�Qe�.1!(��95/>3�;�{@�B	Hg_���9�P��F��#�C4���I5a�������W�%]�[��V��o+�����ױ-�gX 8l+��:��drG�x��v7M��Vw��,U'n?�_�X}���[�8�3�k��h�ŕ69;e�D&�*�wȌD=)JJ7z���؂�Rd}���.�(K1���=}l(���~� �cp�nq���,�۽�W�9]��M��hY��L�yZ�`���AMy�&���꨷�'�L�#�:J�k[�w��̈́"��aʖaC���)�������jo@��
W�nJ� ��k�`5,|3P�&�ܢF�	��eA;a��Vg��7�j��o�%�@�>�']��XU����B����1&J�2�z�-m(�_򂵩p#*?�!�F����F��4����4\Kj2 U��7(c����BL5�n�a�\�Y���A�Z�k�˧o��ޛ u�k-�&��
i��27�3��^S�؋�}u��$p�q��w)����e�J�LX��i�$"I�{-b7�[�`<O�Xн�A�u���s"m��Q���?�Hh1�7�Z�v%�џ<�<h�`�<�f�%�(����h1�%ŭ��;���nB�l`���`�1w�Ì�^}@¦��4�D�����fǢ�ȌL�J�$t��y�gp�N+��G�ew:���B�.������Ӈۛ�� �(�G��8���mC��sυx#>���	N�?�9�#П�WhP>7�g���d�ᔱhc���I�=!4�)��Yڏ��T��L���F>ǌ��������J�~�ԇ�K��k3g�H�;��\B���Y�
���y�9���2P�Y�zp%�$"|(St�c�ދ��s�H7|���.��?�S��P�-#F�����o'P>�0��PA��C�$��8�u��׺bruZ������*�C&>I����8�`��8���R�Y����1K�������0Z�� ��DN�iQ:��Kx8sF[�>������6�|����ӯ�L=�I�M �!�������x�^�H�eX9Q��8�T�T��3z�P�9�r�p�J��,"rƭ��	��3�n{5�@��4�yOWO��*���)�_K!$�w @��X����"���?�K���X�~Jt�O�������D�ls���}^�����g�*ң#P#�\�lG�νz���x�W��%�J��1����H-�V��t�7A�r�J�s�c8!UM=��YUqi��l\�P�"4���Wb$��'���zF�f�œ4}�w����,�1��6�2����S������A��߬��F2���c��aW�y��R~i��<�Е��v�U�:�G��NӘ�f5*�z�\p���o�WҽB�Ji\�O��ʽ֗?������|V�o�p��w����O�f��fb��1����i؛	vu�\��V~l���Q���a�p0S�K��`���E�.˅������IaoٍCd�%���`C\)LEm���K"�Z�F��E%vG���y���:sK���E<�疼0�V]���c��ncOd^�H�( � 9#�I{�@��U�?��l�\�;E�*�(�Ď�+�z�B0H������D�M�A�0<�(q}�h=J*ġKay��M�9Ӊ=�S�7�� ?%��y����w��}�6;! �8��
-���l@K"��X_ �<&�s~��ø����,���x���L�,l"ga�J�C
�	�"*���J�_�F|��:�h>�l�0d�M�D
8w�. A�qI4Rf�� ��S��wt�3��!�|�#8~��Z�a�|L�)�({��v�m����p�j�v���:[��%~��c�Ɋ�ߟ����`�x�~'%ߝ  ���J������*��t<L��cȭISP�3_e�X4��Z$�/�)����G�k6���?���N���k����BC�I�$���oӝ=��?�Z��d�[�r�T_$��?�U���ɸ�Fޱ�eJ�1���㗃9{�.����˯l"Q4X���R����Vgp�f�~�)4�6�I��S�,�������M.I�H���
X����vΨ�E��!
���V�s��!���ڢ@���V�����E��K�A@�p�A�����+������D����؁����y��>�BԺ�k��6.���MDH��G�!�0,`;�j���1�"��M��4��[_u������e�F��<�U�UC��U�G���a�q(x}/���ϗ��5I뱌bݵ9/�"���=�ɋ�?T}��)U���`mx՜��� �|����)������y"�O沺�aa�`\-mհ��}����M��!���B[YX�+��# �7�/)�2_�E;�&�XX�M�!����C��(�k���񀅎g�#G��/tA�d#.�*��t��3j�����H]��>�a�hj�R��
(�_w��?F8*��пs�y6te��g�HlkbuE>��:	��XO2y^J戾1�oF�+7�ܙ�N��6h�0���wB��׈l�>�27�0���ߞ[lѪU�*�����q~�dy�h�D�W!�\�F�}g�A�
C��2�\
������c��76N�Y���_�S��W5����Y�gَ�!!IERv%��n��ڹ�����7�W%�h(�ݭ�J'-�X��.�q�~���~@�;Q���5x�.�dN��]�]�M�`;�\��1��{縙�:w��}=D�h'�!ϐ<S+�̿�P�@�W�UǴ�9�d�g�0CfEHF�mB�E"��wc�5Y���
����Y��Ay��x�e4ك-_|��,8��u������s'��aO��=����6	����"f�~jbv�{��,&I\-%���<����r�_����4GN�yQt���A��L���R��y��O�b�DK�?�[� �f�˥=$`=�^?e�_p���^��pb�s[�u4��݀�_��g�Xo�շt�(��tGs��?��&� <� W|"��3�ps�9�~��S^�r�v*`S�͍����$Vͫ_��>��^�&�7��`�OAᭋ4�3�}H�b�\K��:��E�*Kתr�lf�P�0֌��^�8h;�TD%;��^�)���&w�CMb,_ّ�<�ݸỸK����GV�+j˟SxUY�Lפ=q��5#�C��g}���p��B�h�C�{(��d��ڃ������~=��5��d�~���/K��jC͛��};�����S�絠�i0)���<fmU/�a1@��m�b%+�	JBOQ�W�5�� ,/IP2�K��Bnw��H2�E������i:0����_Wь�a8<���S$0�.or��t���~\Q�mt:� ߩ��aWVkN������-��R}���i@�!�	���l��
�*�y�T�x�K|tRi����-�v ��Q"��Lܨ:�d���	��B�-IcJ���hx~���^�M�(���ա��b,_8����zI��+�M,�:��:9��6��;��hoDC�u�>�uYlJ��ڴN���gV\�b3�	T����'<s���bT�~�UW���$�*���+�y�,*�mLb��_�ѿ=��>�&G}�/!��>	%�K��sq%��*e^=�h=J@{��4P��������,�"g���Bj׷�?��c��č�Q<����%mM	<tZ�����z������xIV����zL(+�|��E�44��h6���6~�Y�AY*s^{�L��͘����F� x� }9̕(���|Ք�׳���	(���U��]`�67-�E�_��1zd�&���&+�,�uX<�<f]Cߛ�����+�0�m�
N���x�~.f����$���?0i����b�×+Z| N_d5.ߦuxOϠKܷ2�?��cS���z�̊E���nms0�tB�3E�8/�.��<��[Y�=��L�pD�A��+�~�tP��=l9�9�-�4�b���(1�J8�M��;LxPY}�.�	�l�5m9�&����ht�� @K�  Ep����i����r?>��D�γ��锆��q���k�T�a��*����o�Ӄ�����n������C��8;&�?�z�Σ�}l|l�=7���@�x}25�n8f��N�3��np��lnݥ�*���/�ݾ׾5��G�c�X�߅y��;E)�m�'u������]�`%�1�4}��r>�*���O1֦�/_�x�j�q}��� #=���Op-\��m���6Z����6���Z��b ��C_z[`�9YX��Q=�A|������kQ���1�5�v2��檐j��`���~����y�fV�I�����<�y65�Ѳ���um䡠y��t_efo�0���_l��[<,k��R���j���sE��xHv�_�u��Ҏ�J��1� D�ꂽǮ�٘�����ͧO���+=�=���qK�� S<�<�Tf?�:`%�% ϔ�5H�5�C`�g߃��p\�������G����d��^U�ɀj��!<AI{�Sa�kmb,%�B6�xYX�2�5�с8��F+T��R��_�B��2���1�z��oy��3W��?�R)!�aZ��9�c�VT2�rς�CĖ	M+���u����9�T>rmE�H�;,^l�h҇��y�a�����N�%��YƏɈ��>��_�K�)< ������Ћ�rp[ނ�)��}4����9;1p�jEq��2M�J[vm�����ǛvH�d$�\n�X_�T����I�e��̦`��J�u�6�y� DOx�po$L�1�g��*Z�z�|���6���+�azψLg8X�,��a,�y�mO����d��-�@!��۸6�}�I��w�Ź�Nc�V��������m���c���J�K�S�rKE�D\�����;f�3�ުڻSR9ξn�y�W��q9���j��~}�v��;���z�7[��m!�[��l"�.��C68һ=�ҦzOK3��6̠)�o��R�����调k�E�{�-����~��\,ok\|�s��o����e
��+�_���V[k���?�;���Y�4�����e'�cݡu�s`����TEl/��QM�`2Y�׫4�F�i�P�� �c����y�o3됻�K���%K������(Ѿ��?1v�ox���餲���` �A�}��v5�b)�{Ȥ�2���t����Y|�1t�J�Y.z�2r�@0�cGVQ@L,�d��\D�0��^ΰ|��|$6��;��X��E�
�r������pW�)��Y����UC!�鲢j����[�k�%�(`�a8��8��6����Cc)��`'h�4��-�I%�7$P}����r ��>W �o�f�>U���P��b#�I=|^�̀zu�ƣ���͍b|��#,�]��
�\,�u\�uMa7�ղc�H�J/��5�����c�������a����z�m���C0	�kk������VT�nՁ2��=�y�����ֵҺ�$���P	l���ͤ��<���+��=�r�Hx�ל�ɩ1~("���R��"N
��j�~�q���0v����ceMO:�5/*ry�.o�%����(�)$���G���8<LO4(�9y�b6��)����0��E��O�*"��(b �Jd�MBF��Ӡ+��9�A��wK�	f̑��9h"�K{KHQ;�o��'�X��@�M�O/P���Ѣ�q͌�qk�H�w;bι��>�u[���5�]Եz(t왵��a5w9Q���5�g6�vCl�V�j�H�^9P:�`m���<����D��-SY��y>;'��&�:Ou�7���Ωf@�����G4=k���T��`,	�,�?�ǲ>8iXU�Uwж���T���Ђ��%�KK
��j���8�Gޭ�$�xs��	��gw���eL#C7�X��I@�G�x�I�ne��Lq?s� UT��^*"�5���d3l��L��U7���:��톦�w6y���<�)��H��y�s׏�0���3nƷ�u�y��ؤ�>t<���<�o�3����#&�I1|�rqǁ��g�	۶H%x���~JiL���O�R��B~��{U�h_���}q�
c�W�߯�8O�p��fbD��3 �A�9L'4�6|�؆���(�#;^��_�	4�Q۬g���*������H8���?補*�.ܩ��$�hO�G�as[sF��	[zx�ǊAy�8�ۋW�x�qhR�ɦ�7��xC�9g�8��z%2��z��:�tn�_&�X�z13{���'D�d���6��(��I��RIB�������Tx�q�*�O�a{��e!�t�x�	��Z�sd��#�ءqc�:����������,0d�D��ȫ�xp���)C�[�QC	��}p/�ϬƝieIY�<(��xx0�����&����<&˥z^$����B*nN��M��Au@��Bq9��`�/��,��	�.�sr�í�v�/�O�/(�_V9,	Η|	��ۘ��o���l����-���i�;?ao�ι�G|��sT���@+u��+g��4���x���=�z�����:�N��X��o<G@��=eVeŴgރ�q��ã����ŀ�a�ڝw��lO��X&sDNi%����ލ��� ^��*!kn��n^�ۯ�gb�lɄ�g�\���E�'�����n�C�<��>���Y�8ڋ�h��^�-�]a�j��E�jhP����3���m�)�'ua'�P�<u�߸΀y��P�9��s_;�.i��@�b��o�I�~��0���}U7r�fWh()zw:�{���V��g��Q��	�����l8gӋ.<#�$�ι-�HT�aV�����ȳe	̝��n	'�aJM��Ѡ�d,��upe�X�l����wu�y[W���	;��-U��n��0
��gEgK
a�x��T�b [����yr�M�y�z'5�i����x>��z��3ǃ�9�I��3<������S,a}D���w��`!�SFg�&�������;�oѴV��_Ug�#��lh�<Ɩ��g������I�l�-*�,�j?��'mX-���u5�'E=��V��[�?6��\�z�4��D�o������2�6��x.^{8��h���^<[�P\��~{�JY�1���K�ƨ`�b���Z�+!�0*B�o�ѧ�C;2^��<�'�TΓ�o<p������)O=�1h����tD�xM���y��S9�b��׮���ĭBp�R��}���X�<g�JR��r֓(+�<L�rQ��6�b�F)�q�D�W�!9��/����L;��*�J(����LG4���Uh`�ZR�%�3&��;�U\����t5adV}L��e�ҁnNCK$��!��|�lO_�d�#kĮ�7.AdIK�q��G��^W��$�V��"�,�W��Z?�/�o=��_6�J8ZK����|���=2�a4=���rq��E!���������uѤp�(v�;f+��K�ށ��u+Ort�[�c�;T����*ʘ��z�&�.Y�q���Da�A\����+jT.�}V�a�[�P8���^�p�c�=�G��5>�cB�rr�����DH[�c�̨�i�ة�0ʵu�#�Q}mZ���^<g�`'�"mB��M��z5a�_E��E+ߌ�!6�1�&��+_������#
�Q~�r4�{��q���@���t���$�4S�#F�Nf�^<�������
�\R͑&�*_=Z��Z�e��o� ��L~��7��8�t��k[U�0AT6:���'�F��yO����N��չ��Z,�����P_U��I������D��ELr\�(t�������Z�x�,"?:���d�T��?��3�Hݵ�S{j������Gk�2��������t�,���4����݌w��&ˎxb/u���Z�G�N�l��2�� I�b�g%4k���wDc��D`y��|�
V̓%���-Ʉ�@���D�j�!�r�F~:�P�[��=y�F��$����.��Vކg��@!"��gL�Q �i�c���ֽ���h�	� ���M�B����R.�<��;Ȩ�7�Wע@�6Sn�p�1��K�;�
��n�(3gњ�ԟ�_�D�o �/�s�62k��Igg�E�V�V�#�.G/����Zی��y�T":4<|_��~���zcw�\i��_1�ݩ�5ǟS-/[d���I��Su�"300�u�P�v{��d݆c�}�Rfe���5���&y��qR}��w�x�q��n}��H�b0F=���!ic�2G��Eδ)sn�0���
2t�7�_8&���a�+�ekrI���`����	�bk8^����1�5�*~��Gwƭ���"v����𞏤��r;e ލ,l��'M�E|q�ɫ_ߏB�w\k�;c���7Aj=K�J@1�n����X���|�����Lrp�$
,)�V/�����M�i-�����x���eŁ���D��y�L2s]�U�D�xs$���q�$Շ�5��T�3�0��8�v����,��;F$�9.3����$1.�w[�����/t��R�Bl�[If &ΞΟ����	�c�ėtۘY�L�����>��-�-
�&^b��d�\8N���5�����0*N%:�C�;��ɚدT8\��E���8�n���'Q��N�X^D��^���[��.k��e��Oy�}`'�ͪS����?hk�g7𿞘����ǡ]#��jʀoP���s�o��/B�x3(����#<|]����&: ��0���;���p�Ԗ?��RG���r�	`���QO'�S̹?&�Sg�f��ɳW�~������g%f��y�ӂ���F H�œ;�e>�6?�׺/>�/>l��g���"?����4�_/rϒj1���W:N{��=^`+%�#6��ZeXlxV64EB    c291    2010�'��c_�W���M1[�E�ZT-V��2���Gu���3Qh�^c�I5}д�N�R}�9{��B�Pe8���?����� �mD��3����b��T��7�7�Q����y?�W�~b
w�j+� �F���2N�ʥ��I1{�����VD����:���&�fQ����K_�<��GF��VæOV�~f�#Ѿ-� �!L=��;��C����@��R8?�V�U���������\>�Zzk��o��oI���_;����CV7a�W���q��~�J�a-�ҨِDɼ����}��ڬ�\ �yk�ީH,�ʐ�7a���2(�QQ��Tt>j�>��A9��)�8��I���mk?J����!�P�z���ƽ|ʿb6|��W���C��^��Ru��ŴX
�D��0V��jc���T:�>��]�����P|}��j6��|s�>á�=��L֞���ui���!��n�m��|���ۍ%bO[.nBR��FPs��s$�� MY�̾�¿ڐ�?$"���(�J���K#�E4�J���2��&�υ�>���q�T#�c=��F��h�o�%�+�g`R��S�X�³%�i��/1WS����j��!p�$�Dk�>�u���:*<�e�>[�������*���ȏ�}�&����%ҥZH���G^�Z<��פ(�
��ڬR]_;�N��>6���H��꫹Z���xŚC�u�tn�ú�^��z�	��q` i��i��Ě���'<h�s4�?���٣��ڛ-�/ s�Ŏ�2;hTxmi��	�c��p�\��w�����x��HHoM?I2|�n80��4�uE�G/��^E�h��h��m�7i�,�@rR_���	���7�+�1�WN]v�,�T�2qY����J�&p��ΰ�ʏ���*b�}���C��t��ƭ��]{�N1E�'s�y��U�m�a�[�c�x���%��L��P�����2���)�A���9m{�j-�����AUԴfG����@ڜ.���O�:oʞ�f��L���ȄF���(=�]_�6�į;�n֜��؎O�J�'��"'����3)��dR��7PiE��C������(����K1��=@���i�_Hy߀MH��i���{��k�^t�x_%+_�gk��c����6d��Ƕ��;y�)E��������u�A-�B��1�}�L��f��V4�3��N
c|�,�`���D����Ǌ߄R��C��hV��*�G�!��R�O���w��GI�39���A��e�A/ x�/]\�y
�/�1 �ѵ���=mVc}	LRP�P�a�^~Z��'R�G�5���뙘L���ZGb�P
�v�*���m�T��=�!]G�H0Lg�ȫ;$H�����WJ�@�j[٦לE�$)�J!.2s�@�����d��l��R���bQX�Z�U��V��I�����A� ;4[��Rt7�[�U�DI+ �W���C[�>U����6��A��|�;5�do�ms�I�$i\�������T�H�jsi�������KȬ��,"����X�Yid~�U���%���|D���<�3ףTd(y"��`�.m��?�f�B�LxU�'��?���o%����C��.U���,i?�^N�g��*�3��&���8�����gbW�5�k��>��7)2g������up��^\��B��>ۤN�hG�P��0��М�1L�ߧh�rzz�h���փ��N
B��=���{��]IfBF#�w������̤�o͜���~�m�Ux�H�a�����ly�/�4/�}/�a���O`���5�C���`�nE.��zg�]�+��V��B<�\�]�1��
𞄊�"W���t�7���h�ïv��?UV�����=��j6�S�Xi�A��s`7A��c�]�Q^�MJ���#�M9�'m�4]òO.���G`Ł��ճ�kd���S,��@y�b�o�)�r��v�>����h%��R�̎=���P��8�ׁv��l�� �ћ >�?��C�^{>�w=�M?��������,�uj�	�~�O]��!JtLҐ5oM����"��o[�����0�p���'�~g��;��x��$�a��u�V�T��j^��������әzzދ?�BuI �'u<�}N�ƅ��b�ǁ�	\��*�2ze����.E=��W�T�3�����{��#e1p���_0"�����33Ϳ��X���z�V@�'��sM�_L�-� ������#O�Fe[�1m��!���9�<�����m~��+�i��"A��{�p�Q�=��)˻]7.��! �p�}�=?��N��"��HGY
��u�:P�km��X
�fF��K�u���U�E��+c�nV]'Y����d�7�A'��U X�Oa�{[�>�y�JY���p|�6�
?V"���x���@3��n�mI2���_���>�'�F]�V�0��m@�(^���5N"DE�\���l�z���(�js���g��-�o�лG���S�R�<�����"��6i��*�8�J�(
s��Q���ZrS1��AA3�g�Ԟ�ޫ��tf���v~���4u��u
�x��#���W S�]���)M�~�dZ�
�ԉ1�#O/$�u�[]���f��_re)�y��&T f������[��{�	�)�|$����n�T	���1t��V��&ݏ��xg����At��qn
^�f�����x�&��鏄]x!�3`�� O��M���R����/�=����w�k�j��w�=Id��~޲]�_9�6n��b~�S����<+��%���=�=W��2�g�/�j'˹�hOa�+@*l�H���7��a&��{[���,T�k�	i�������y���B6؛\x�%�LD'�zE@������G:��%P>��<8w)�)�._1�\(��?Զ�3W��@��wk�<�W55����\��ݤL��c��U��P+�f��).ׄ 1'�\�qu��?
�lW ���2qU��J�����tͿ��4lzL`S)3��m1��0	W
W$J���C�V�'3�6[#�!]�GCS���ȅ<�O�����.���_ZN��t`	�O���t��ш�4,�B(�Y.]A��J|����;�F��(_O�G`E����h�0{R��h�Mhq�@Zg/�0jPN%TQ�S�wBÀ��tߣ�h�ޢ�r�:߼4f�����"KN�͟K�����q�0��"v�:��̴��P	$yͱӱfKY\�� �;��܃�-�V��z6zx�P[��S����\�Պ�DA��R�z_Vus%28��>��<��*+Px�#�?���D���_�p��eH�2���j���&5�A.�[��ذ+;����s]Mb!B�K�6,N�G��{�FF|�n�舧�~��ċ൮2�q�����/�;�B�z��j㲖������L���@���"�\.�Z��UǷ5*�������!cSY;$�@�,h}��v��t�:n(d��;�����we�](�����s�u�9��:z�:�ʛ$��È�J�?pLrr����o��|��g��Z���S�׀�ђ~o��_T��nYt�;��РN'���9.�z�B[�����; r�Eb9�Z|��c�����d$˙OԒL���%�)]X`pD�@�  ^���Z%��Z���ം�٭��T烱�`3���sJ`��s�w�����x�n�c�~����x\���X�YN<��Ә/���Źz�Ŕ^�U)N(;8�^,, �i=���z\��?C�"�ΪԳX���ϡ7+���"ݚ�1VM?x�������əqt�*2�5���A�wf� fb�r b�-�]x���<!k�=�Q΂���6��/Oحc���Pf����ïJU�۷(��s��4��M��P=sOտ����2Xq'��_H���h�%%�.�<ڭ�H7m�.�9�>����� :���p����OSŭҨ��t�/5ޮ�c�,$C��a���7HD%4g�c���
�GspU�È�~��a�|�g����脁����^P ��۔
8�}��=C֤=�'��ڴM/ k���3s�X�G���U�i�#Z�!�������qh ]�2�Ƅ����A�{���k�K�ag�g�� ;3�w5S�ө:�"9
	�<2�G�`c���)�t!�4��(�.�]��E �"ʕX���x�#�t
�X�Yz[:%�9Z��9jO�#*��x�a:;�!�F����C!��ȿfgCÅ�n��Cj�fZ�0��VMb�� ����^YM�� $��w����?g�jpM�:Ͽ!jl*,�7�R��[R�O����<�M��A[��C�����eG��Pғ��Y�pb�����K��;[߷l��M���4Y��:4Q��L �ޯ�t�-(U^[�
�=-�\Eӳ^�]o��./7:�8���2�
 +2��Ӿ�j��(,���j�)�|����y���=�m��N.j��[�{i($ή?Co*�`���M�#g��5;�[���WA��������_�D�-+�Gk ��w�O�c�Gǉ��mh �#3�I���Щ�k�:p^���������ɰpei�|����DA�����"���r�M_�DQ?־���bM�>1nOj{��6�C��������FM�F'�~RR�T$�c��l_����/�2�w,���L��� ���@8o����O���JTQ:,�O`�FX�Md�߉�����/7�
߯��k���"Tϼ`(�7{o��-����P�cBɑq�O�'��%��}����Z��E64�w���ո,|M�J�hK�1�H�O��L�v`�}�P<��j�k �	��s9�ߐ%;mm��R�暔��n*%�%}�����vg��x�|�E��8��@���|!
qt���[djlw X#.�;f�u��C��?�GH��M�?C��9��`I��kV��X�Vh�@��Z0�e��ʐE��>��Kp�P2祪�v�9����k�S%��U�����}]e�Gլ��:����)9��u�����4�積�S(=�m���CQ��h�~�M^���{< ^�S���hDT*9�o�6���!-B���Q�&�=0�*G�m�^A\eo��L@Ҿ�]abS\�v��Wc�O�e�Fެ�}��X��3p3���b8ɋ�&g%>xx}ƹ�9��c�G��J3q�4F9t|�{�b��N����f����Z�|�:��ɮ��~|���^I�����Vʊ�� �ǉ,�LE}cǯG���6���Q���N�3P���� _�0��:��^��z���G[iٱ��yt	�a�Pq��/�l��[�w�IW����
�L;%�1�vJ���#�錖�����p��겉jn4���@�B�ms\���E�G�,cչR�`���'��7�$�˂�	vm_�a�R�U�dt�\�/���I�2��������%�$h��������C����� ��J~���tG�L��H�#�E�1n�"��k���`_\���H�i[HY�~92�8`-K��͎����T4eme$%�ƙ`��F-U&J��lK���"�S�+�]_�9�St7���g{����d�Mʪ1�+�`~�nA�(ge��r�A���+���s��=
e���f�V����i����5��G�AWղ�lO���ZPL�23.���h[Ќ���텣���kw�e�S���vm��f+�
���M�9�D��7�B������_��߸�
�v��n�:.�T��x|wM�L�%&��e�$��K㿔�ã��Nnr���ba@��gnf]�o��-;��0�TWM`�l���������Ly���ˁ�x��	�Ju�p�At���
�gȧ}چ�RM�Lv�!��sܧ#dz�럸�G��1q�7-"T~C�V�L���[��i�����_�-�Q1�)������ [c@D~�q(J��Ӹ��鴊(���1a;�������ѩ@.)'��U��6�b�ȔFo#���E7�p��8���7`�c,t�6]�+�t�Q����U�7�uR��s
�jW��<���Ʀ+.�k���0�Fl��.;� ���elFy�N���N�?y�|��4Š�P��Kx/D�f��S	�"�{W��xP��Ô�i�m-�Q�u#9J������V�
��r�R.7#&�gs�m����L{�(�Z��~/��2���T�ˠ�m�r�K9+��jRcx8c���D��m���9���]���l�~����d�g}ف��bD�c�{�ī���4��Mj=|�i�
�}�� �b���H�AX�*�f��c\�	U��)4���Ư|4���{�E���ܸJ{b}&X��D�{�[������W���P�@��J��r�z��5��VaE�e;ժg����
�)x���r�{k䖚����N}��ڊRV7��hS<��>��>�(u�����?�ܘ�h�ʏ�c x\-~���mpw�4�ܱ�1�\���C�*`˳�'�����2¥�ͪ��3��윔˫r][�v<���N\2��׍�D��}�Q�|���X .P�C��2�0���g���YCu�)��PF9I�ʥ�R�0�	�שc'��g�(�2b�\Aw�7\�X@U5ka�w��
#����	t פ��VA8K�ذO[�%��'4�W���	�qO6"X�l�b�阔�uxm�>�����4N�	�z�*�{�c�{��>�H��cBԾ�`C(��-ě�V�k�00_ �a-�29y����o���y�w��$�g�5�����$.��3��s�{�7G5ʵ���qZ�:؉9!�b�0��'hMA2M���R �DRG� N�~�
A��{�����.[i�����*?T���u���
�5`�Yi�Z��(*1kO���o�]$��~v-���J�"k�R������J�uP�%�r�w�樓��N�xJ�*�F99�dq6ۇ������*H�=���E�u��̂�	,^���w	X�#t%$-�\�%�6�t�i�W:X�lh�<��g^w
�0�^	�g��+�VSG�2�cP<�SFXi�Ȅ �.�߫��q���H&f��І�v�Fy��(�b��o4��&������QE0%���_��� �5lk�%?��/����{Sݜ`-����l�H��++�'���|�zL̖�	
���\f��F�ź��vѯ�&ɲoܦO����nwI�^X��!�ϩ��� M����%@"��L�|
,X��f&�{9b��=˨�2<����q�s 6�8���φ�^�Ӹ4}�>*b�[�,�^��� `��ɰP���V���垴�{TP�*=������F�t�D�݉^�D�Éz�
�>��P�e]zu�x95ۏ$ca��T����ƁR23,�r<�؀����Q�u�r1�P�`�Yɂ����Pg/m�U�w�;�x7��č6�����%��I��*�Iƾ��+�����]�N��S~d�:ob��ȅ�,yHx��򠃊*:�y�;Faȴ�,�g˘�����@$P������S���_$���1�io����%�y���iuQ���i�f����f���m\��%M8���X:C�E�q���4n�r |I�( �G��<'�}�`�Z~*��MG���G4T ׻k�� (a��(�Jƀkc/_2Tg���-)B;�g�g�5��y�:�5I��,~V8ؠI��kR��9t@%����3��M�.�qF�٨7�j�e��E��K^�5�=D97��C׀�����/A.�q��_�8St�q���[y���y��� �n^�����zآ���^��6�M��U�+C}����_�6W�c
�6�����jO������-V,
��6^}	iez�uŀwu���1��Z:-T��.�c�r��v���3�7V�'ه|���,���?���h�hT���7�h��d~�x(��|<�[�E1G64�8���HA.�%�7�sܷ�.�BG�A���[c��^[��J�j��0O#'�k%�k�F3��_���TR�Z;󇀮�����I �ltr`~N�7f��%u(mgn�\�Zz�Y�x�g�Բ�a���I��J/