XlxV64EB    fa00    30a0B�6�9��G���V*�U�2"3��y$�f�	�h�ggzvY�>B���r�gU
�\	=A��'҆Y����5,Z�ty�b��Q�
����x,IvT���ҋ�R�&�ھ��8�S��}G�Sz�v��S�C��;�kdu%,�����Ѱɒ.�Ը�b����K�AOÏ��;�x��*{H�ӥ ��o�{��]g��=^p�ѕ������H��D��lj\��\(u߁q�����W0��{�'���_@C�8�0�cSS:�0�
�B0K�1��3)Pi#nG$)� |y�ʬi�i�N����$�rb�>������z���Y5 ��a܊d%r ^�[�y�R�q�(Ԝ�)z�ө�:T�.���~l���c�(W��~��*Y�\��A"эOq��n��zU��Zu�e�:K�Բ�[p3�^����]SS��j��!98d3*)?���+�4т� y���]����៿��3�����翇�Ƿ�!�"�W���R�׺����g�D�# KDFPW7��s�yw�U�mP����W����y�߲��I;@�p$�D��m�c|<T�Բ�̫~\��ȅź�����^���IFײ��40"�f�K�|�X�o�!����H�9�Q{̪%gZr]�=�k��4`�9�&	y�H����<���ڌNưqL�L�@.I��F���w60&�hW��z>�p�է5]�'��� �8ߟ���|�ڜ�'U�x8�y���:2j7��U0.11Z�	>�-�{��rǪ�	Q�`�Kc^H�G�A�Y�����ثпp�{�܇����h�j�[�q�(.�͎g�Do!�E�fo�.}�r���AD\��x5K���֑1�˃O�
F��(#��gj�.�a#���[0�{�%�$Bʥ���\C�i�Gu]����
 ���������>P����/=�GX�vC־)�E�<�ZIڧNN e�;�	M��0��|f?a�'�]���s��n��Dd'̍]r8|GR��o�S��}�xN:��3c$,�P7�cUх>9�{Z�Eb�؞!=JV-{���Lx ���� |�
U�|8פ;�v�����牼���͆��/<�$M��<��z�3�v�^���!Qb_%�e���1��pw<*�+q��WR	`��ʧl�d�E�Rĵ�~&�3P�L�{�@��zK��^��U�v�������Vs#+�R#@GM�0ش;�ZP��o�[7��ӕ��<w�pg���y�Y�d�q�"����M�v^�&g����	okOw����2TU����L�.(,�I&D�D�3xv|(����6��铈�:x}R�H��ŏ0?$��$�����hQ�ÿ���N,��t�V��x��zcR��Oz�qq&!2$�I?�!+�AX�v�m��8���gI�p�����o+�v$<�J���H}�ߓ3J<����<Xt	�G�zt���V��^$H� �S�K5�v�[��������\�Ѳ\����EkJ����NnbT�}����>��� wr���K�}�g������Y#�L*4Z�6�M|���l������9l�}����i��V�Ǎ9Ӑo~�%�4�M7����Q�I�b�C��P�G�Gi�==i�VF������o�z��jW�Y_��C�f;4TU���꯹O��e�$����h�ڪ���j�&��&�bq�Hz�\ -�%洿duhC����	q~D����eG�#�@��3��z���Kk׽S����/��o���`�dC�3_���BI�zЧ��cP��C���J��<��J3!�Ɍ_����%����7�<1�ʠ��bu�&�����������,�/ބ"��&�	�eb���Fm��&��)��ӹ�~+M���1��l�Ş�|��5�-�fv���UV_�������Ċ��q?��dvz@�'@�-�M�a���?��k!#�i����9�^�Yc.��Aȗ��lǅ03&	ғN��l1r]B���-t
�P�������=/��~���r���/ .��Jx��F'(v���SK��ɝ�9=זqݦt��2�a���k�/��5�$2P�\�V���w�=߮r��s:�Fs&ef��L��R��i�{�o6;j��~�O-�'�ŸCM�رY�# � �PM �ߎ�*�#_d�u���%4��Ӛ�7���#��65��)�
�=.,��B]�䜇��j���_�^�A��VD@�&{�}��"e����owmQ�N��/��/T�~Q�R""���(��Vu��"�|*&���4F�q3��&&�����!U�ٝ7�lTet(��>Hqd��ծa.j�q�y����߮�x9�;Z����})�]�BkB�>eUȏ��l���NopU���4���諧`�����<���{�{!\�+����c�s����&�\q]�/�m[OG����T`�2���ڈ�N�ү���?e�w�1$��̨B�NIe{Èm��2����-�>ŅF��N���"��Hi���rP{�%����A"� SE�@�:�x؈@� s�Y%��;#����|���b�S(�H�0a��iW����U���u-'6���{V�Ŋ,�B�O���y3ӝH>m�J߲�U�׏��n�_��"]�6��t�l��a����<Qgv���I��6ˠ)���K�CZ�_%�8�\|�F�u*{�ˍ�}�!� ��]$0�ރ�"N��9�)_#�{XʯH�$C=��u�H8���i��_ć�H��������Y�2��jy~.\�~�e�3�ܙ~(�8w!�����\��> s|��OPlt�m��r�z�i�W�KO�s`E��V�p�&�|
r��vw�~n�������R�!g�7�{(Q�rx3O엵V��S=��q��[�^�"�0��fZ;m��$v$�\U��t�j�����2�t]�[��Y֦yJ"��i�BMAX��"Nٵ�U�8\�He�	�udL���=� ����dq-�H0v�����&�R1�9A����ez�L��x���Hv(��,c[2yf��ێ���ED1G�|k��+��*�k����	�s�Z�r��������# ���ƢG~l6;�3�l#��*|�AͰͥ�[P��Qj9��_.-�KPv��0����੿x��
��f��"_x���MwN-�e��<��׳�Ŋ��`��g!����(��XF��̄���V���;3͈'�4@cŚ?6�������������v�$Ou�6�6(汗�Q�r�<�O,үb�
`�%u$�f,N���A�������khJ�r�\w�W#��Ф�x��P�t�N:Ƹp|\/���`�+��KV�	���G�W�ႵO��B�8�}T���8���$��S�q��氵W�x���4�#np�)o=�h�|.�;�v�;�v`r�W�D���ie�j�oE+F��&gC	£��OT�n���Ǆj`�;P'Ɉh<t2)���K
!<ʙ�pR�Q��V1�E���
��i��bi�6x��!=x ���kRTþBp�a�P#5��D�?��kZ�Z;��N�+ކ��r)�8�T�*Y���g�~*;��;�/x_�<�0�ig��1%��;#϶��E�v\!�4���̾���NF�-1����M���C���C�/B�:��e{'�'r���)v��?C<��M���c,�"��#�{W�>��m�w�I��U������i�c��D�D+�AT�]�Y[��&������-�R�&z�_��G�!�e?O�u+�Cׇ�9˟�ԍD�"�#���u"�-i��� i��^�!k_��VK} �+yB�4����#a�"�;	d�L9/r [k,Iͨ���hu��Y�B��P�?L�}��q�ȫ0_	��_#'��.M$��C�3��z���;�܉��sx��J�☏��1������T�u����<Kd�K5� �:B�~�ʇܲ�d��[A��Ď��Kو4U[D���}��)�����`şZ���,J]Bx [���� '5�Є���b��Ύ���%��@�Ȑ0����=�9�yN?|X���[b�D��QB�����XwK./<�j��j K�Ҩ϶�^��xg�p(>ʬ�<WBi�b�bo;�t�i8�붊�FׂC�06�ل���Q�qZ3�f�����^+�x����߲H�#���K#կCˑ0��)_���o�s������U���|V�yx���"7����T�y�r�ϐ�����/�ް�����9Θ��0�[��� S�� �䌼h<Z19u:��_[����YI���%�9ß!H�ew�,Dq.��A���6%�o��'���5 ��Q��`���2D�2�������Ɣ��������jXQ�:l3�_\X	m�=�_,�up����������/^<{/Rj��7����iU�!.ÌG�c�����1��T�n#�\�t��Kw����y=��e���X�pR��k0Ux�Ki��C��3�LB0ﻛ������(N�7l��P��k��T7�,���}FEtN�*�ά���ޚ��@��@�ӔZ=U/�X���"G_��_��r3�+��p�2g6M����|�lRY����3-j�4|�5�܎3�u�������E2�ǲ
�'L��RH��Z��"�s�BY;�x��z��7�t	(�:�Z2�K$c�<��~)V�� z����oF�E����dm�/��ΰ�������UNw�-���;�bɢ�z�imM�q�~�������Sk����v��P��,V�9Ǌn��j�d��j��� Ϸ�a��y`9�t�[�[/5�pn<A<�_ޛ��VI���.�Bf q�v����i}$��>��2�	̀��~�����\��'��M��m"��:�P��t��t�JfJ��u���l,v/����v�nw���}��2"C 
�j7|r{%�b����'7� �MZ��G3��g�0@��fºA���
yÑ0}y����֞��K�2�j!���}����5��Y��Ӕݧ��̻�hwWg�qf�
a���di	����d�����k�d���Y���� pV~6$�g��Uhp\���R�[�FQV�.�H=��>���ʸWz�1\�p�Ok/T��S,��]�+s&]���/t=�ԓJ���o���U��x.f��`���C�>�@��:z<켳�P t9'd�&����ޣ/��%[1���?���t�$±��:��X��W�Ɉ;���w���V�V?�yDڜ5����'9��e�a�#�ӣ�*?�E��HL7ND�{�},������;�������dh&��	D�Ơ ��u�L�ҽ��9ɟ�*��F+�)�\��q�B�c�z�U_u{�5r�S���'�[Y��0�!��?�u�=6h�L/���kY5�77�i[�t�	H������(%n�E��<#58Ѥ�yb��vM��\D)�S��[b�Q����_H�C
9���҂�}�3y�S��ӰZ�m⻨�jEI��E��$ިA���9{I'nڽ��+�爽�gr��?�༂
Ob�o�i��v̤ȏ��3 K~*��l�5���ꈼwO�3��@Ƌ���T�	�s.Sū�=+�}|T�g"�d�M��|5\5��3�
��R[ߥi�C|�0��J#N�ػ��ST �䅸?b
Q���K��O[���,��Dy'GfIi\1n��0���o�"3��}"U'�="����7'��*��?�^O:�kI�L�Jڽ5&LY,*�4�����8yP����F c�"NdO��
����:#(�skd�oZC��v��R��i�9�L�-���1�,:��M� ^�L�����~��!M#O�4$)q�6)��v��V3!/$�L�ּ1&x�4�rO�����b'[�,Dq6/�O�9QJ���㎤�|,x�	?�u�ք�W��_�s��)W'̪(��ߧ����U{�|��0n (�����]oD�I�,-����L�%G��uY� 1o֍,ߣŕ��sB��X��ï���R]�n�M��/y�zQ�@��j�R���u���~Â.���c �cO@���R�� ԇDv�?-H���?|�YlDu������s#�˞E���<��G�
��(����<a��l��2x�f�is��ρ��f��ur�<�^1焀.�ŝJ,�P�ᖙ�f	3GM( d|>q�ʫ�u0Q�+S}[�˗)�E��v�C]�6������>�C��[�)�]i�}����,���F#= ��U���eF��9�Ҝ��E4��ˢ#a��{M��g!����F�0��U-�f�.��n�2A��.Ŋ0h���N�M���
��\1�w:]r�?������2J[��eX[�!��]�b������Is�bS�O�Sj�I��	x��������
;CWo��O�gJ��3B//IG<OOv���|�����:��q���IZVa���P�)}&)J�ʛ���"����.�?�`�7�P�O����W����ʨn�Z&p�}�51r� Ro敿�	�[�B��z����_IGv�%T%�ܓ:��d���-�:�9�ͭ��)7��/�	�J��+�C��t+bC*�Tݙ�gU�����$?维P��q�ĔӘv�R~�� �?j{Q�?X�d�����2PL��#�Hg���R�̬����*mmK�P��ڮ�"V��o��
�"���WnN�@��p{�Sb�	o��\ȍ�� ��J�h��(� �7{�] ��E`(>�a���s�H���aFk$�D�}-��l-6��Q�[���5^��.0{���ЃV�v��:i�TʗB�>P�ˍ��=f�t�,��)t#t;�;�|a����[��0x�JF���ׇf=�����h����|�CF��w���6��=��ǎ���5و�ޝ���"J�~��}�P/1 c+�b����x�:�)s�~N�}4M�AЧr�2j�E[�W�r7�]�����E������<��'�+{R��2�� ǡ�3�D��C(	=�5:�i�s��������d�X�K/�5!����=�u���?KU��Rܰ%�4�_����xmf���f�,rQ�@�G�hl�M������z��)Z4L�iX%�J��g�����^�;jq�4q[\��j�w9��!��U��m��[h���X,� |���OG?�BeVQm��_��(�ʌ�&1�� �����cqnM�#Ɓg��+���J�r�~;�~|�w�93);�X&7�^.��%6�	�=��Y�]ǒ�*rJ�ş<7CR�ҩŮT��[S��� �Ƭ�p@EиS���fX���`$�?�m�21���N�u	z�n)�甾���5��	�j`e �<Ta�%�!�,p�ՇTrh�.��n�=�j����0s{P�S*�3�|�PY�A����PPkI7?Ԥ�2|ûlO��b�&8=NQ�>4/�@Ċ o����JJ��x��)�3(�r�T�ĊG��My�7$���0��q�9���=�͛Nl0�Y_�gGt�z�upG�.r{��гR����	 �:�bOY�^���?rp9��թ��%U�����$ä��5�d>!6��΂�ϚDk��/9����˟@����%���w�֤�^�U��1���q��R27�i_�@3��9�4C�Ҏ8��B,����J)&�Ӝ���6~�6�;	S���/
�i�Xe��
b��Q���EQ6h��*�,^@A�ɕ�͔|�_b �Wk7��� �1wb�C�l�Д����_\�_
2o��c�._zI��d�h�#�vt%��VHُ�ߚ��D-�y�]�	��#��T��]�,.Y��YR/F�,��L��W	a�6痼E�O��Ъ Z���yB_��v�UZ�5�B͡��m���C���Ȩ^Bw(O0����.�Ә3B�g��,���k�<�� �ʾ:D��?�>�Y_F�]Hz��F*F�9g{m�v�Rܛ�Jj7l���A��r����7�� Xc�����؅'g(�k�:�NoS5�\i��hѰs4RC�ә������z�Ŵv�@�a�� ��hw��$�fTx��(w^�):�Ej�M��@1X{~���M�'�{�������]�V�Z�jS���n9�B�b��dG⮜,�@�\�\��]��*�R��k�o�\4H)A���f�]m�c��)Z��2²����BZ�����7S?�0�t/�`E��2�@bn�1s3u���D�������f�,�hסe��GyJ���m�/Y�2��-d�Ҵ�ݗ�jH�x9&���j���fQ�Ie��k���kk������� M�lr�[��*�5g�������k�Vw�iX>n��,����$�=7����s�_N�T��m���/x�G1^w��w�?��f2���97@����`�����|R�2h���s49��\R�%eo�ӱ�ʼ�$E_(������,ٯFN��LF��mk8����ڛ�e�Zȏ${j�?r�	3�b���?�Ll�آj�,8�sc�h�@v�}�S��&����󊫉�$��"՜�E1����Nׂ�J������3 �s~����X)%��������m�o @�/�%y�q.t�yS
�O���W�+�ޭH�ˈEQǾ��V�O�����Oy���|��:����U�ֆ�{�1�(��$������G�ĮM���0���ݰ��p���9,��Y�{o�- o��s����􂢱���}~ ,�Cy"��rn�����b��Л?n�w���@��Sg7���� %�$��%��U��Ф`A���Q�'6��޶P��M(����	t^�Y�d�=�R1��N䢞"�;2�"�|���6 ��p-3 6b���eW��d�����a��@�жT����=�='}�f������X�g0m��k��[�.+$�C����J��&�S4�l��s��aU��WX�@kΣ�i�/L�S Go>��w�&} |��}&�i�,X��P���f �F��KEb���A�=h�B��BcCU.\�� G��\�$��n��Gؔ(ȁǴ��tM��0Ƌ���t�"�����OVU�B�gQ��*�C�)>[�FZp��!GB�O���]���崲U���l��I�2�{�*��I��q��
��z�s5F�g\XZ c�L {��2���K�u�n��%��&��v�&+O�4OQI�@��\pڦi��E�x�└�*wK�zbы%�B<vīl�>�"F��bo�Ky/)�����	�9�rQY�$�w�۾�� J�[�q�5��兆~�* !W� �æk$�2��}�����T�GVI����[������1��OQ�?�.�J��7S���z�!.���!�6�q�sͼ���1���%3�V��_�_8^*��tm�w���TjqƗ����W�e���sL�L,K�[������>[v�(:�6�0������E���X��8�X|�P��������U�� ��p-�kLdn���h����O�?����_ �8U�R'�1&q�s���U%F�E��׌t�4�$�6��T~w�7[��w�D?�U.*�4��ߐc
�l��2�`��wh�a5͌c:9�u�,��g�jRh�%h�+�9���04��g���FX&�D��P��m���G����L�og�g
5clW�$1�h~���w��eR{�)�;�`�vy�U�~�V5�L'H�?�O�I��Eȕ��'ׯs!�pq���ʦ��;�!ݎ�x�B0��k�����]�|lk��k2R�@���Q�`͞0� &a��_�B*��0��x[k�(�Y�D�WmcY$�x,<�񏢷��$���(��k�}���*�f� k��_�Ď�+.G���#�+��v6Ț��\;s�������{�\v��=�2;��6?�yE.M"g[E�Ԃb~@����~��<��Wk����ߺ���NU�$�ݧ�}�� q�skUb�-eq���ǵ2s~7֤V�� �����+�c���]Ԛ����3���u����zA�ǌdDð�.s�J3�Jq��� Q��[��r�)@�Q�gA�"���'�^k����\{d�h�ܭ�#�q�8Q�����Le�w*e9Q`c��̭ �s9�cXM�]u4�)i5�L��L�Va��C(Mv���UNmB�x�Э���_�{t�~j;f݂��Kf�Ҝ(�ò5q� 1�I�6U�b���ߞ7 zhq�Gz�i�[��S�,K��k*�^��@������o'-�S����Ukx�#ٜ�� &-�����J)��,���9��������G�k�&6��E�V����y n�5`"��EM�&��a`?.�E��>y�І�X�7�4�lJ���ZŌ��l�z�oX)8��w1�%zT�j~�5�C���'4���q찯nJ�ec:��	��E�V�h���-T#�[P���^��o*f:Q���sN$����|���V���7��JM#�~��"ZBV}iG�����^g��iH�ZƹH��s�dn��)����-[�a�Dg�Ya��c�=%�;@0�m��gu��sWh���
��<�W��'Noſ�2���Ձ�	-�0W=z{"���^�\^#����װJ� �`�N?�)Ks�d�<X�����^B�����Ӱ(�&Y���>kJ(=�R%D�Qpyե,
��������sO�/|��+��L�8"�4y�j��Gm�p�gH��� sv�=��C�Gq�l�Fް��j�m�9����L��� ���)���R
�����Όs��ids��/�����Ǌ�\��םY�7(6�.oeA7�փRS��G�L(��k^:v�ׯ���͔kr�dIQ�������6�C�3��fVd�Z�R��&5�b|ۚ�V��W��-^g&�}df2&P�عG�3g��JBs,�l���.�l�s'�[u<�xn*��+!6Q� 5͔�� ��0�V1�T@g�vg��'hi0Y���ߛ�b�hp,��$K�/�.��w�����Y�(����	/0�.�h?��w�����"��<`��|�&��:{c;�'���6�Hr�!�$[�v$^3,�#���I�z�
�����T�Ib�����IگKE�[?l�{��ѝTщ��%�%O��BPK����nC $������R���	�����\ �#�O.�6J�r���C��Y{e�"��m�ѹO�	C�5�->B��N���h��Q��{�b�����/�@�>�ޅ�6���]�����o�H�r��>�y��6��;aMY��w��QcTo�ҥeD��O�:�K��������kH�̝�x��f|V�FR!�v*Gr~DEw�v�F�H�$�i��Ugl&�eMY٫�"m���h�4��*Z�6h�#��l>�h]�Q\b\��n�d��x���Q9�y�^�8e��jyh蘙��f^"��A%����#�۾9�N��f�C�F4���B���ǁ*굂��薢��ɸXy}>��g�B9+�g	��E���]�+@a�~�����$�(6a���ꥺsp+�mQ�=Ht���-��i"B볼	������\ƨ�����H�tk��-b�r齚������c�瓝]��g�w�Hm�px~{�\:�:�%�I��Jm���&�x�S$v�g��Gj8=�X�#䟍p�+���i ��<��릚%Ķ��Jy�<�`�d�ܢ�(ly4��(��h	�x#�t��)���~��+���ы	�^�Xp�u���/\�0����g!���[��K�e��}+��*\_��6�#9ٺُ�L��R(IJ�˰�3�;������r�U9ɳh����;��w��6�Ra ۹p�¾\հe�\�F1o����X���U�J�\Ժt^�D��.�_���l�75��2�`l�e������~�$6�6[����U������ᎂr������U�Q�|��\P˸/�@E$��xMqo��v��Y__��[���U�\"��T�Un=�4qq�\�̖WHyu�`����	B����ѳ��Zot����20��XH�� �U;�2������n��bl�,(����5��T�~/��7on�n�sCV,wJW�ѡ��m���X�(��M��m�V���7'�֭�1oK -"b��V��ed��'�󤜓�Q����e�Aa�f��J!˸3J���P�&�\�--�-�r!�5�,���؛0�b�˱���AH~[U��~f���:������T��Y5,��b�b�2�ծ�IAҳ�*�Yc�v#��"�s �ۿ
����P.�Y�2~)�s����X�XlxV64EB    fa00    2ba0ݷ'4TrE�-�L��K�b�e�Q��J�]��/)�ڜ����Q�%�:'��/��_ϑ�ԗ���?3�+�K�1�D�n��`��:���Ӫ���ߪ���Fv�����p��$�W+��ҝ�l�2nƕ���T/�L�=�q�P�]JcW�|]h��-��=��m
naG��53��&�uhλĲyX��fʰ~�����m�6�t1�.l�%7̭������H]j5mZ���g�&�v�5T�:$���<Biψ�� ��|����S�����=z��1�	�Ǡ���U���V�L��_xe��ƎQ�����yȇM�oz�]���RCҜ�0�����"������Td8�� ���<FG���a4p
{ӮDxoe[;�>10!��Xzn@8 �B�^"ÿ{%�kd�3�o��̤�q�\U�܎6����A*�6��p�Lw��c,@�d�߭�>j��`'��}��M��W>9Ԝ� iَ96�D6/7\�'A���]�|�8*:ݿU����HT#���` �.��9�v+��b }��O�{ّ�  �';����B8��xb����ST������NK����-�$C��
���#��.[as��
S��Pڶ�I��kOƃ��Z�[�Me���{���Ȫ�+�m��&��2�w�*�R<x�8b��3�M�Q+�Y��
��xJű�	�x�6% �����F�8#�L��5��
���d�a���@]=C�ࠨT'��k�	�6PnO��5F�}�D/�V��f]�R$ Rp�!t����q6�E�f��䥪���8�q�4���62:��?F��sKib^��}���du��B�8�z
�V���vPxT��z�	�W)�s5�y�a�:�g��/����`�:�W�J�	z>h�?�Y��?�P�faѶ���N�%U��K�V�<�fO;���Z�%C�I�喨L�'Y]����>7�����i�ot �G9�
���((�o�l��;ՠ�Ľ��J�]��~���@�mH�z/���'>�^K�|��n,�g��%�2]�M���IU��;p�|8Mݺ������Q�əq����Ы:�N"b1���<o��7g�_�h�lc޳�y���R�h�yt�R��]b� �t��1�:����dH~&�&�S�1�:y��(���Nd37��\��<�Vf�y5`�4$�	�C�`����|l1 ֶ�h~Ƿ�m"[���t���E8��Ǎ����Ygq�?A�� wHV�:$��Zw͵k�!h��≄�6���n3PAF�}Ft1� ^�L����&��e� _��h�{�*���*ƊGZ����'�%v^i�6��ID-v��Tx�'ɀ~�<n9��z��nj�j9^�e�l&�G]zY���-����2ZmzV����AE�|�� �pwSa����vA�"؂��氾��1���������ق��B��NI�Z:"2=Y嵬���j�mԋ�vA<��l���fS��}�U����8��GH Blx"X)[�UcMI�!���vAw*z��L4�?�5�1r����n?:�E�)��A�,>6�����y?g#D�(��!{�{��i��Ǳ���(hEI��(��g�9��=�H��؞&dH�q�Pt��G\�4R58f(1�^�(�S��r� �k�x���`DU߹��G�5�wu�\��{�1n�b�����x�[~����*�Q��D"���e���r�IqL8P�C!Y���]h�+���)fܔ���1�bƍ|�{x�05���X�s���3bu��m�m�{�0(P+�~52�q�<j���j��|!y�3��%@Fp^wD��zt`3�ynl�8~h�I�n��V=�I��Q����	��n�T~{�#��^ 13�Pur��!�KB�a���'�h�γ��2`Ϻ���0�3�s�Uތ�����޲�A?p4��9����)��NN��B\���_�X���v+��_8��=.l>=����_�3sb]}^�H^�΀����1��BH1�{���=���MW���r��w��nu�����l�<���a&�� �cH���^�$6 D֨��n
��;�1>��\dM�1�����§����i�^�RJ#uL�K���={�V����z�Ŧӡ���b��p:�<�f7U�(� ���ߛá[�KW��UG�4-;�Ϥ0(r�{i`�������3�&�5%Z@C�H�eAx��~�<&�V�ŊË�x盋-��)��������&��:�NyoU��т����Q������[�s�������k�ϓv�.�В?�u�`��`C��^�o_�'B��J���/=
�x�ZvQ�:n�Rr�u�G�=-�t� �7���=.W��y���jSh������&blZ?�}���+?ǵ��D��[|v7x�q/�xlC�����[���i����rFźȣ4k	����Ol1�������z�1=��zK+��%M�Q]�����i�[N��zg��� ����R!��9 /��nh|&HNs-�Kj�a��%"C�����9:��
	���~Uw�h�i����(؂��д���}���jq밍t�Ϋ�&�����5a�J��`:.p��%���`9@ڄ��&��X�}&���O�J����V�-�PϠj�j��]Bn��=Qk�FU�@����������g]���i%�B�`����Q�{�����xTU�#��#8Y����~���H��a������tSMo��~����%�|���.�a��ku��S�O������2��ѥ�� �.h������a�"';k��[���*�W�e�H��nPs
,tҎ���ό
ш�Y�)�D���k�gyy���^��Z�5�K߰Y���S:a�*	b/�|ul��B����a�%�����r�1�N��M2���v�0�<��ӕ�^���3S�@�;�zq�@�6w�U�.n+sa'z����'#��|z�
�,b�Hc\ϴ��f�ƻ�aęF\��ꟊ\4Nv^u��|��ݴ����H�v�R�����8J��8K���>�`�j��}N��˕B�������L�r��J�	��� �H���xyڞ}'�
���B#����*�D�Ӱs�}z[w�D�dࠛ.�/�E]7dB6V��.U���qx.u)h�No�����w���E���m���_CLM�
ʎ�.�����:�<'�H7����X�Y����c��l����t�ł6�{�P%(����?P�5i�kV#]S9{il�z	S�r�� 9�R��1�?���"���}i�͑Ґ�o][!í��6
S^76���U"���^�T�~��n�2*�@N{%��@�2�sQ��G�4��H�[����|W5Qs�9�(��>Pd}��t�Q��d@J���G7:a��[�'��M��yy�m0Y=�zUx�T0�Z�(B��-�*�Z�.�ϵp=/��uU���1	��-�� 8(2>*���{���l��V�RA��Ɂe�aV�l��!�� ھ\���z��<����2��$/1�A�����1��*����	7�>�]��F�[��lH��e�_g=z~�E��Vv��R=sQΚ*����a�IY������qeFB�'�� ��橧������&�S���L׊H���Lk�x8�ۼ�b���R ~�4��rҗA�d���;��~w�N�Ĳ
q�b���C(�X�5-�L�o��As��SX>(�}�.pRd��F#�PoY݋�m�}�4�0]��1o����7'��(5q�#��D��44��T<�P�{�ZIԳk��7lZI���ǃ�i�'?�,6�����n�c���"��PB8o�d��B޻4�B��U�m��Qx���0��m�C<���Z�r��D��p�A����g7ܛ�em��&�Hډ�8�#M�������ד�'�s�@)�!zu놄I�A�85���3D')��'�R��0��ًr�3���T�����yBw��r0�Gv��3x���4�4m2��	8P2���� ���l�ס�{�9�(���v7����.��+R�	7��h�R��.V������@6��lvH���"%q?x���w��bL����X�Q�V���IDg`�+��Dt�*:<Kpw�h��x��{���.�r��g��DAZB�G����?����kY~霬�(�I���ub �����-�Csi.����ސ�_�I�Oe��k}:���&p�����5�~sL ,ͭ)O�z}�#�,b'�S̎��C�-��6�ש��^a��&�a�4.Z�~�*C��"�0j,��[�q�aB$�zV�0 " k�rܑ:����*��B]DCPߔ�t�i�q�K��}�^�@`W�ڲM��TFxCo9}��s�:��'�KxT��}��b��U��\�ߥ��?T�Hb��u_��g�a~]c
,���dWZ@F���<�ܹ�GZ����8��dg23�<F�����e�(�Ԗ��>�n��;�{��;�8Ӗ��[���9�<gt��7�O�q�=�G��@�0�%Y�[ݞ�����^)f�B}�G�Z�/�ԇ����f8��x�E�qf|�}�{I���h;�be$i�0���0Pki�BO�ǗW@���}�s�T?Sc��)�jq�kն�݊6ѣe��n��d���"���pǓW6�z����"_ǥzy�
�F-��I�*�:��|�<��4�J�K��*���"���^�����Q�_�� I�r�ďC!��p�/�nE�(�/�@��3�eJ����׏e}�@� a�m�I�H�	��r ��E��i��#˼�s�W94��9����5kF�>������ D��CqV���-#��BT�&�����h�l|�{�)�
H#3��8,�������W�6���?@Q>�������O�s��R�{8�nF@�Dy���Ma��\v3P���!)B};W��ߜ��@(�A��'_���V_i0��ќ��&��J�}�r�E�L�s����ള􁉪غ#`n,�Ac��t��4c�8?�!!�n�`�=�.-�5{�{����u�)k���Q�P��(��Zϳ�����W��Ǳ�V�`�z����/�)-���,�{��_WY��w+m��r��ؔzO�/}��V`?�hMig�3ڏg��mctGqV
֓x5Ld<M��X�W�Y�0ex}#�Y�i
3�]���o�:�;���,��z�O泻"Ջ�PL4 ����꺕?���_����U��c��}I����V! ��N�V ׹w`���E�wy���^�t,t����5�d�����;R^�QvQ[
~pu݆�@��) ���e�� ���2�ZN�i*�`���|��2���NL�����	�ҏN/>U �����2z�������#�_F�99�֎rQ"��R�!E��}����D����څ����Y=�D+��Ԩ�!����R`����V\"w����'*./���\*v�6��a��̽KW�@mY�W����l߶��e�o��8�����X�"Aq�� ���|�Ҏ��U��Q�Q>�೵@�o���R�MW��=#l�� Cxmz��2�DR,5�o|y�5C������'���|�n����*L��:���[)�d�m ��<��E�h=]�Uz�QP@��'!n,$]C� W�D�Nd��=Y�RE��S��N��B�2n�$0���"%�^�Hc��Z��!�٪HC�k;M�����f�7���V��6�zwp�lze�;[J}:��ĺ3]"�a�+7����1X��������ʬe���4�v�_�6�IVh�&�h���ɨ|/1�/�_L�M����}*���ƻ��|�V�?�u�x5�����l5��qW�7C��D�����[�	���y,7p�|�ї+)	�K��G�œ`̛\F�E��!?/�*N�7r�≊��gJ�LH\|�F�����!$sq�#�N�:��G1���+J��G�Iw��������b������n�Ռ"�+���J��lRv�LU�[����Fe�^X9�W�I�df��\�9�q ��{�.�������c!���ȼ\[������l�%��	@s熶�̻t�?0��z^�	P˿0��f6�;�",������N�-(g�R�rz�*M{>��9{)�9mcG�>{@=y�{3�|\����計t<}�C��Bw��)XЮ�s��D#zm*��<�:ja��+Dz��o᳉�fp�8ǩٚd�"����E�kǧ�#�?�QD��Cu�����)��7-�&�;G<7(ś�;��ߺ�8�|��,�������)[]-(h5xC��Q� ��'ۛ�_ך� ���	�c�+@���f�<3.X�1gW.�0%]M:m=(�)iH�{\�[!6����D٭��^���^ʦ���o��ާ:4)�H���V����2�[���͟��@�]��F�=0
����B�'E��d��ݕ��*�df��-=y]A?т�b|�RAo�9��{��݃l	��u�jn��||�k!�V�z���b��odV�����h'Z�@SV�8�%�ߴ��H=�E��F���
x�;$V"��
߁GX�1�IY�M]Z����׉��Ȳ�+r�MHt3�T����t�)�0]����IU�A=�
����Ʈ���:���?�-��ʛ��?k5k�S�֊BR�ryJP���H��-��7a2����?�6h��K?�*�����]LZy��9�s�?{3w!No7E4ȑ�TwCt_��P�{_4�'���zkڮp=�a��e�(h�è!JE�sq��$3��V����8Hz<�](�=�� �UR�!r9dɓ�B�e�t���m1����?с�&( ���Zl����:đL�<�e�o�_�4G�+����
M*i+G#^Q�̯��.��������.k�dܰ9��{ƴ�>�����f�J6���l��.�&�@Q)��|�vqX&�ѣH�i�}g.k�HQ�x@(,ܰ#~��:Ѯ�~�C�������֌j2%C:��B�:�����3ꜰ���&pT}X}�Z�W�G������Zkd$�Q����ÔCҨ��7�[
ǮYE����Aѵ� �@z��5f��=�l�bt!���,%�sE�\��#�Q�������]x1����wx���lChMKk�.ב�XaW'���E�.�� �xq�;f�0Ͼ$�O5,�c������T��"�	���}���U��h���z��֬�̲� �x� ���K���:S�a�.�/ْʰk����30�����9d�E��ǐ4zgRM�"r\�>�)��򩶧1��j��3fEuV!4_��%�)$�F'B����RL�9���Ç�3Y���\r�7h1��ݦ���,Ix���XgF�v�y�#��B�W�1汌��I�L2�:s���[����m�塁�F%�押(j� �!���|�Q^�Ui�ϵn�F��~E;�����'�l��(HY%7i��š}���6��G���ʹE�(?=�u�|��/7��7���9#��v�Cs�t���L?0��[
�f�����M���J{� ���3�P�\��6����6u���)sln�lx���4�!������;�A0\��$)���
gH:�#����y�@�\P���=Uj6S1��蠵mۚK�$�1~�\�9�C;sv��X1��c�/�������@Ǡ,��H�GG��]͠{�3�cQ=4���B����4�wU=$�+�G�����]%@5�״U��^W�#Գ�P�\R4����hFA���5�[��*�:T9�ۻr�r&r kiR��es'�$ Պ��_���w���o�[��省K��M$�x����t�'L���S�����U��x�P@~+��,ySTȸ�1���*FV	 m���ʣ���Q��E��>K-���z�B������ eҨ�а`1��?��������[M|=G���?*�p��n/8���-]�Y�<��D1c��f�o_��b�*��k��
ӧ5	�g��"�w��J9�`�^N�p�X�1�%Y��.���M���ܺ��W��2j�����+�������t��ۃ�˜�Vym�V�z9�������?���(}A�H3�HD�o0�f����׶�/0/�B1��K@D��m}�Lyv���l���\�f�l�S��i~aw�a�`̐��R:m���]tD�fM�e5�uD��Rx�������u���Y�<��$�O�m�(z��N}H/����g��T���G���h~�O�cfv])Ws}��}�\��Q�Q6Q}>�^W�/&zk�M	�=P��*���mE
F|�]���v����0�z-��>�(R�w ��ۊ{V�c������@���vW5a�@�K�o��\�Eq
��~��24�Z�s'���1̌lW �*EOqvt��OIXE�R(�l�J���7� ��ԕ��;ζ�Z�k�F7!��{a��E�_�GM�����`n^qB���9Kyb��o:Cz��Q��)w�Q=�r�{"�����&J�<h�]��2MU� ���G�r�7N�~�`��#{�<8��
0���M2�<�A����:����d�YC;��H,,M��"E��ɾ�=��+vD]��[;��ek/�9�B���8��m�sr�� uN,q4������Fj�g��;� M�+g[�m� ��=K�m���R����m��qKk7����_��솙}0=��TWM�44���o�͸���h�O��>~�������W׊�D3��ޙ���]ɐ�\z,u��G�nv-���U�+6�,��y[�ʨ�"k�10f���B���~2)�^��{J���2Q����\�0#\�e_�
�4� hfІi�u��E;�Q��M�\����<��j.0��2�Y4ػ�5�^ɼ Y��T=�*����|B'�J� �h�1�y(j�WE��
͍]����hx�b��N�qR�1;&2��kΆ�����A(O�)U���G���Y(�0E ����c�#f
���,5�H�ƹ=�ѵn����Q��rٸaQaQ����s�41��T~�����i�ɬ5 ����a!2YQ�6(B���béz��o�g��$��2)�����	O���M`���v���yƈ�ȅ��Y:���c�\Β���]E�`�2l)��d����Y�ǐ�hǟ1�i�:�����+�
�͚�o�a����|$˿�꤬��rð�HRW�#gP�AL��E�/��mq��P��sp>;v��P�DS�Yl��0��/�&X� ��0Ѕ��
ʄՖ(3�s��/�"w"�c7��|bs���=h��O[; Tx�R����Շ�!ô(��&uO�z,
�kӡ�����m�|��Z��ݩ!O|����#��s.����L��ʝ��'戅{�$��2�7Li��J,����Z�T\ F����9�r���I�����$V� �%29"HC�	�:�F��[@����	غ��BS��1A����y#i�������/���n�?�|��b0���91��`&3]�G	��1[�S�o"��}Vb¡xΈ�P�X���#���y�����]r�Ʊ�_�4O8z�8M��pĢ$?㘠��cA��N��젤� ©��,��#z��+|n�`����U?��	�XAh	P9�$[G0g�'�������s�����0�>�s{Qp���8�F�4��.4,޸Y�F-9�;��m��F�����l��_�5<REZq��&V\@�d�y��e��dލ5f�p�e���v2N�����f�8��b�%,�=b�n�~�����7ɝ�A�iro αrH�Z�����pm�Y�� �����g>���t����� �|c�dh�#�돚�ms�o&���f�E"��Ϛ�W)1p���\zMK��-��|�FF���εu�]�@͆���䛨QO�o}ΐ���Z�ӄ�vn��I���-�Z�7ܾ[�	T+��*�B*��b�B�Ƌ*�F%�1A�̞��Vus�Z�k	c�;���)�����d�%Cn�7!���;	AmKmQU_���}:��v����l���yc	�kn�� �ye7!l��IxM��xu�/�C���Ǆ϶�>�M�v�VO8�f�\YPFʊ.��/�,r\���@���q���X���Q��7�谞=�'��SvS�T���N "�A�0�">�_�0ic�\���$���B��&�\bBMњҖ�hT�.n����U���x� ��R�/SC�����Ih���Y1-ݛ�~�W�-,�E ��&��B�ҏ���-m*�����	�/���,�p|��ʣ{����0�T:\̼�?�x��U�����I�TWsL�%w5�[ҍ���{x5i���m��c�O8bԱQ��������7�ᐻ�C\V��N~YoF��Q��������W�	��y�_�x>ݑ;�,�1�@;��?���������U�H�ſ^�]��K٬�u�����&������.�=H�,� ���g�r�)�f�k�����1	�y?�*�t+T��քH�x4ƚ&17�pV�"]��7��rܣ�?�8)�����lR�"ˢ�JQ+��c��ۮ3���ɻFp��h�i��3&�)oXi��q��	��,��k阩���q:40��n����Y��羸����B��&/�����-m@��Kܡ6��I�Y���N��� |�N
Z��'%�#BR���9-}�+ �₷�`��
�4�.]��,� +��� ��U�m�^-DD��w�]���֗��ܧ��x냤Y�Y��e�p!��w-Fk��UC������ �C�}�o�i�N�n�Ly�T�3�}�P4�$�g� '�k�O5}T��:�/���*-�zE=���j�m��>cNcp�Ȥ#�(u�c1wHP�ϵlˮ�1��#��+H�(�-�ti;�u7|�%XlxV64EB    fa00    2710k5";s��"6f�7��G�*���l�ؚk�5(��+��7���S6b���[i_5�F�p?S��G*�,f�i��>I���ݤݣt�g�ߛkO�=,wm���\93iJ+�5�C�<�P�� ]��Rl���x���'��e��UK�]0H��Mss���+����d���skLh������ rE�\��4� �6�2qmj��	!���?�Ȕ�����\bo{o,�u�&���+#Is8준9�'~�<O�e���M\9M���H���ĹQ(�Om����x�g�K�qؘo[	M����������S�L�F��7�"l��Q������R1Zh&�6�O�����oeZ(ID�����;e����a���CZ������aoj/Sq�7�j��=S�查��1�l�x�������H7�D�T�F`�?jjB��h�vR���Ӟ�I����E�������7�ܙ?f���"�`J����M��~.�
��>T�J8�]FI��,�ے��H�ؕrR�W�����c"Y�f�JP97z��rvm~��']+�l*�fi�H��b�:�8W��I:kQ��q�$�P��P5~��l=x�,"j{��=�de:�p�7M�(���s�.���I�7g����n��:��$/�D�r����r}�ҕ`�q�X)���,7��@Ks��0Y�?AwfF����,Ŕl�Zc�3i8��D��{���{��ՠ���F`j����ض���ʨ��^0��.|�K�n@�T"�����/��{��ה$�)`?�/Qp���z
+��ЖG�3r���:k����`�X�Iv���jh��Ն��	p7�%�C�ص�^`�a����lF���4r��[Z�V6�(�/��P��˚���ۚ�;9d�΂��A�n��\�El6�S=kc����ѹf	���F ��z�R�;���!iP��cǔ��jw禧 ��w.�c�Ӑ�ʹ.��M쨻�f�?&Èi�sG4K��(��f]�	�C!������zM��V���-��[�X?��׾�����zA9xXՙQڠn����|~���G�Zצ��.�@<B_o�.��!mh)Cɚ䖯�G���N��R�����EsQZ����&�����ĹA3�e9���Q=���|�����a�J�ԝ�����"�d��OV�B�_��[C��,hlk�����8Q(�$���]U�?�셙��+�d��d���B&��3C+��E,��%�\ڿ�MU�ǎ�.e��n`��1�7Fh����'���^��ѱG���E�W����ސ����R���
���/�g�����ЂW��F�=�:U{��lM�x���c�[��@=}�r��A��
��M�o�{��6�^m=�=��@��d�)�u,����	Θ�"y���KI�2x��@���=�a�??�%hŉn*��
�^�q���S�f����t;��56߸v��`�>�hi\���Av����-���5�$XUףm[��ژ�０M����>ly9�Iv�^ ���^m[�I��=.;���'֚�7]���z,�ƅ�H�WY^o��,������ظ��X��jJ�}���MOo!{����f.!�<�_9|l�Ppb�uʊ*y�\�Q�Q�����Gp���� կ��g�-!o�*���b\�q���j��c$7oDnي���ʒ�ךv��ݗ���|1��:i�9^9�T�Dt��r	�pJr漕��C��$-y��l7
����-�!j0�bז6��@���~���P��T*nڵ����©�}��:��A=��9��_9ѕAU�HW$-Ph��h��������L��p�T���_m~��\C)P��F�d�t.� ;#���w�oUO��#�wF-ȟ�P`Prܟ!��z�6+%ƍ1
��38���b��rօ��F��8O&�I54�~XH�q���!�����uM�Fzev��\ x�+�77֌
Bot�U֘i�;ǊE�	i��8��]�ʠ�]�ZF���l�+�`__�׊�<���N\��p���<D^��1%#^�e]R��Ոv	~"�*�OK�g�+��:m�d�6�T@�{����.��5Ր��jcS;��cr�-��_b�p�=Z$�c#�r�}��C�D�Cʓ�����f6��������N�7�z�bj���Ͽ�0�|4��]�JsF��1���[�8|�D����9i����Iw{�������Z�Z�����&����QƘ��Ȣ�0��K>#�~_&W��uu�D!�?�&�浔0L��%�ޡ��HE���5�12�P���a�@�. ���Aag��kQ��Vl���_c����E��y���}`0�����5ya�,��GM�yy�B����A$F�۩�����k��`U7`}{�.^������y����=I�B+�����0z�W(e������#��L%�P�l�<\�F�{��~OZh�(�T�=W�y��,��Ai������4�p���dȕ�e��%0���~h���T��}ZX���\�u�FB��@����y��귃flY�&{�k���=G�B��� ���ɢ�u�me+�7�j��t�R?X��y7��ȸ�c����je�cZ2]�o��1��]ȵO���J���WXҚ4�����'�oc�K<��=,��-l )�%6��`��4#�2��t�� ��m�����#J��ׯ����=LQ�"X(��{��{�	����'�]_^ uKC���,�\��̅���6qf��ُ}�\%}�0CnL����(G�j���J�r�`ޣJ�����8cP�G�0�P��$͖htՊ ��������Y����̬�s{㹙=z@A�dJ����QRȖ�c��17�T�Qgu���t�>����!��(��T		@�#K|m��k�WY/U	�/\D �I����q^�5;�B���*�e�룰�r~��ϭk������B�I������gڭ?�qBfy1D,ؚ����ν/+����k:qf��N�S�8v#�I"Y�m�\&�^�)���H!�jSj�x��=�~��������Jڦ��zl����h�rIz�-���qH[dRT6G�B��كv�K[�4ۓ���o�G�*	��~���>����y]%���e{�Q;��gE���[l!><mVS2`	KĘ�*ؽ�`�σ_��Y�a5u��O�?��Y�^����5�I�W�B0I���Tq�G_y�
7J��eO��w�ڻ+�6^��_���q�Zq���%��R�ّ����wf��ˉ1/)��<0�,QT�t�.=Z����Oǣ������ܺoN���@/�a��L��"i\s)�ԠF������1���q֘%��e�� ,έRK\��~BVfqБ��e�~��卼 }��J 2B?�'ǀ�������T*���Rx8�o�/4����D��Y���EL�T��#�א��0�}�?�o��3s6]�poE6V�u@�ӏ��Y��[����6��e)pF��%pF������B���@��Q����0���At�#"1SK�Ӹ��GfJT'b�MFVi��y^�������'�N͎��ED��u���5MQ:[�q�-�[~K�����{�Z�nNoqm"���?�M�GW�|>���(���n/�LJ5�u�j5��)2�{�?󵳲����;@/�_�d1B|���X�(@:��	�b6x���,ο�	��(+�b�*��B���Q�� d�1� ޚb`�P]|��r�[��bAk�,4\�0��BhI1�1d~p+����Ei�?2��	�ݚ2�Z%���v�
��j�t�Z4�˯���[r�n ��eP{_�Fcm]���3�{[�i�	Ep�|�Ԕ_N�	d�rsoP|�gB�<��U@Þ�����F����*�S-Z�(J���i	3�_����O>q05��x�����?m����C�3�>�8���p��#���<�ޓ琢s�,)�n�^�tP%���s�P�ػV�b|l.'d�#�͞�(I
��(t��C���i��t��Ӳ�]�%�'�i���1d��Q.wr�,�G�)�L���r�QI#M_��-KH�#�j�=O1�C���@s��,�'M���w�����������3�:���C�0�;[q�A;� O�d�����2F��p�\`}<ǹF�r�dO���\>�%�>}C�0Y�a�v�b��#/Lc���6���V�)e�|���%B��qy���,�y�h镽�<���/�O�a׺����hӟ�{�����̌��#<��c���K�F��;��
ܘ}�~腣}{�4"L������p���o�HC��o�����~ip�+۶RA��E&*c^���-]qI+ן�~�O�׋�=���qƠ%z��ţӓ�c��`:Ce-4vi>�7
�xdM��406M��&U0�!��Y���붌���,��JB����?�k�������\�'m&=ཊ�����㷉8�@�� �s�J+���K���i�,*Z
�b���}��Y\������H���u�~��[�ȩ~���!"k�3|ڜu|�a��t*لw�{�������C���-+�c;�,b�C��7_��_<u �J�&L,l��^���qL|d�ly��l�o�M�U�-Cy��?�[ڀ^
܆ZH!6%c�Y� C%�PE�,��}*qP>��!W�A�� Q�vq&_l�������w!z��Bp�a(z �;l1�-��Vj+`��ȏL}�m���J5ߩ)�ؑ��V�nzJ>y`�L8&{�-o��DuU3�H&7�����H�E�2]l%l{0K���asʲ�U�c]b��C+����������&ݗ�����U��lrÄY�0.]�Ls}3�j���y�f����ۿE�7O��3̔X���V��Xl�|���k�r��ҧ����x,��%q�����s�L�C��7�{�$d��p��	Y�����$Y�0Z��x�'�
��'�����tp�la�$>��IZS".Dn�bt60�B�3P�ڕ?��k�R�t�4Ț//vP׷�d�-���{�����0����#GK�6��b.�R����;�Z=ly�����a,2�R+$��J��~!1�JP)4¥Ro.��ρ��1��R���� F8c"�]t(���t4�XƷK�8�N�&<^򟬢
�u��k	��� �ؖ:�b��Ĳ�)�"�zJ�*��QlE��tL�}G/������aNn"0�ɧ3��cGwk'c�~����Ք�7��2�AibT�]q���?Ԍ�n=�5܍� �堯-v]���܇⒐�b�+E&�"|'v��T����ЈW���#�w!2O.��&�Z`��mX��4�G�p�U�j�)P�,�ҍ[��K��ֈ��ˮ��X��RV��˶���P���uiu�1�!��"D#�� [�,X�'�A8���!?z��l������Q�tl{�Cǘ�V�!v���h�J���}>�z9(;�lrv�~n�D]�:�@�X�/��>U m��Y������=�̑�35Ccڏ�i�A&M�Y{]#[\���7�}l�,S첥�Z�!Tq<�*���cTU�.A$��ݠf���4���ibz5K�e��W/7*����cEC`�j�n��`��}u%����T�
��Y���AEkr��jm��U��ʐ��!f��j�U����!u�zl8��� D�3esĞ�@��b�P��N��d� t' S�@��Q��Ҵ5v�wd�>�Q� ������z᮲�VH�� ��S�g�����~��J��K�(�(�{"(#��&���u���O�|�������Y:��_�1+�-+l�\�u�t�$��_��9ՎL�׈�N��o�L���_��:J�Q��-JE�m���"k��(ȭJ����~dhY��J�y��u wI��P�8�(�	e�տ=5������R��A�{��z��ǃjT���]2R#w�KJ(��l�Z����RV���F0�N�.�(֟!��^U �D��@����\,l
��'�M0�G�=n��n�p�P���Ϯ�n];g#G7��*���>�y�y��;�	��$@="�.U/#W-i���w6gF��dN��A�E��gɇK��&>�=֟��P�\�ڠ }�=�'����h�Bش�.����� ���Q|�L�^�`e�B.��'�2F���fS]G��^J��f>#��A�'6j��E 8&��h�i��)C�y��3�ɷ�.޶�f�b�7���M��h�y�����x���uw����`�Q�e�[�+> b��p�f!J��w��������P��V���ZcT����!��;gLh<W��}8��q.���"�{Mʣ����.�,�m�S��0�ӵa�z*|sB���ˤ2�
�°�]�7j�t�(ЧP�}ĕ�o!��^���;f�o���̓�+���A�-w������b���c�����j��Oc(�Y�Z�]1P� ����l�a-j4�-M1����$�]qC�bxcM?BZWv�1<�=:���n��Ý�oRs^��@� zl5�]-�AE�	 r��a(:^�?��a_b�����G�ɭR��u�ϼ) �;��0�u�]0�x�#O&�0�g�5$S)�P��g����\��f��߽U���+t��l-ֈ?�at���ϱ�c):v�R��<�y�e\H!��>��7,FJ"IR.�ƛaꠛg���<��6ǆ`3\)�͇������H$��}چpݯX��`��&�D�x�G�C�\N��m�Ȭy�ޮ�ZA�F]4.��E����V��id\�Zg��M V�aY�|�V&��r�0��=�?�C�ₜ$�e�o���Pq~>ۃ�����$xA���y@S��ٵ����q�$:��W�'��	Sau xǕ��r[:;�0�9B���B��u�C��3��am9�c�}�� ��Aζ, �@#�W�xI��'kx��J�`~^���/k���9,a�B�'�d�:vЙ=G:��"���9�\sz.����*y:zMAu7�@m,I|=L��xS�	T�>��!_{W�w�$���G1̥G!���wt�$E�@��;�Pnˉ�Kt�iFQ&�)yQ��؝�_�hT��.�8�1�m2��ԭ��O89����iױ	r.��s�
����nSF��iq�tZ���	7���8�w$ 	�T�����s�K_0��u[ViF�yєJ*�㇅�M2R| 3�|���J��e;�*�����GΌ�x���	`ٲw����}H������n�n��e�wx2W>��=���;���jGK�ĺM����\'���f�Y��r8{H��T��_@a�9jcC�޾c,�)5��D�a�$8*��H�{S�}-~6aS���2~+cu�iJ�XB~A�K�l'�<?I�P�u W
�.L&���L���C��%�f��3�&x~�i����Y1��M"@XBE��\O5��j�Þw�XJ[D?���m7��;o0���u�m��r���r�7'���wM_�1���}��yB�u_����g��:��FF�����&;��c��.�Ȧw��/����ż�47���cD � �����!^	4�n�
��gn���Ή�������:�d��_+T<N�A�ܛՖBn�sd�8A�*�����Tz?r���3�����MwU5�Ⱦ��81
���=͔Y�@���hޭs�4w��S�\��Hـy��eZ6�Sl�e,^o�$ȋ�N��嘵b�&��t�P��q�X�X�w0�$|_h/X��V�հWs���}{�ɩ50zW��U�~ ��2�"b�OY�_j$T����:��9B�Ȅ�L����s���y��zy2���G�,���U�/��s��>n3h};�������j!�ֱ����Z�G�Vlw���P��R�e-ˢ�w �%s�ov�tv3� ̆.<jA�`�o��;�RO'����a�*��S)�cڤ���3�A����|�b�Nά��&�p\�@�ϰ)����hW��vV摘�-IxƸ����?b@��0���yy����7h�򗝒x�Ix�ab����(���J>xSX��eo$̘�AA&��}hbo����{��-[�"
��S]G����"j��3*�gR�pU|���hC8��W�,ӫVz�:�D�f���,�����;<���Qj����pUS����[O�<c����L[Ҁ/KY�_%ԏ,�\�ś���g��(/���Uc��ݯ�o�����E�t9��5�R��6,�W�6�cr:��X�Y��%p�{Dօw�thF�2ExR����d-Gf��#D���6 �#0$�^��WY/~���w&U�vW: �6&2�%:�B��c<�h����Aٛr�49�G(�b2���hԕ\���Zj|�#�o�c������#p?X�Y��2�F�A�F!WFs����P2��$�?m�֢.�#��T�I�*f���P�`�8�:��=��c,i2�q�P�ʖ�yom�w�D�m+��􆝋d��)����R)�����	�O��p��i�Ne�P�[�} Y�sz�a�>m��GL�{�o+���"N�Z��Q��6FaA�2��������O�/x��F�☍-�a{]Al�Zl`w\�SW�p�UQ_m��ކR�<�:5>����vI��)/�*l��U���ҫ��| ��|�����S��1a;�u�Mc���I�r�/EC��/J8���愭:>���vڢ�l���+x|*Ũ�z���*up:�ݞ����~;d�B����@g��� Ajp`��͠�8�`����� ��:%I����ĺS�s���"��h,�y���j�JwF}�J��>�{L1f�qD*�z�h���	Xc�έF;���q�k#��L�3]�V�~Fұ���\���6^� {bz1��n��TC0G��~E��d� ����'<�%��]���΅��s8 w҈ؙk�~(���N�(������� �遅��lkv¹�|��tly�����DS���9��)��y~�<�-����.0�L�pꯖ��7�Wr(#nZ*�������L���O����U0ɘ�Q	�W���״H�Ǽ�*�tZ%8Y�����_i><�0*9����f�� ���燼�V3�zp����&��K���R/!.�b����p��t@g�'�pWm2z�X��U 詄��-��rqs�P�2��y)Հ�i#����	<����h$��rK��$�f����N��ndX�-Cv`#26?A�<+^�z{��m��R��!(�i�����xڒ�8~��~��*<�p�e��r� �pv]\vp�*ۃ�h�n���ӓ�!��,�v֨���\>��M�Jk+�P�VHsl�-��1���#
�z��PǶ��aw�УYXI�k���/�A8����cf�u$N�E2�Ii��Dj(�x�x�;�e=������m�>a$ց���~�H$,p�����+��z����XK�Hh+�V�Y�*�D{~���n�x�^Fٽ��{v��� 3�=U�<ұ����<:*��/�,��80V}��jqv���N����AG?�o�tU��a�oK�w�1V|�	��{ ��&B���v��L���&O)I�lF|���N�<:��u6��$�r�N4������s�����S����كWS�sk��ӭ��>0�kRq3�3����i��-�P��"�?5�&l�>Y!$'""�ڇL=�0�9��D(�sq2P�ԢA��]HK���VS������n�n�x��t���G�ឹ�Q�q~.|:�\&^E*�S�ņ����?kM ��� ѐ�D�L~��AQ�� �O�
��FǤ*[]������HV5��З:S��~�'�XlxV64EB    fa00    2430٣��W_֜,J��^���(���r����'�f,�G�O������|���������B��R ��,��N�bX��P���Zp��{�໼YZ��(ͬbE�K�w����v#O����T�B�|,����,���2_�6��Z]�K:s�Q��a�M,�XQ����M#/5>�����K~Ԣ�itAwsm�o�5�4p9]vh?}�'����=9� N�b�E��\@��pJ�:�>��KrG]_�ﰅ��s�"ex�?�,<�G����,r��v�8h���8�:����57:��~�R�c�Ա�Bqh�O3���j"b5�҄+j�s�H�u���Xa|�P]�Ϣ��f-�Mi���Ơ���`d��	������C���%���3K�������|�3��"N��xu;1p-'��כ�[��	��R��1AE��UWx��AP`���y�a+�n,y��GSoK����0�Z�>���Xv��4Js~+����0�8����Wŭ��t�i�.����u�S���C?0�<G���-�[;Iyf�-��@V@�C럂���b,�Ͳ��e�X�,^X�,��Q%'�O��:����"�7!͖�6r�F���V��F�ə��0�	_#^��yN���u�س�p^�d �4���&����<B�B}�\�L.��A9hn���M��I�0�+�S~�5���X�q8��#�?w��^�c�k��i�����
�ů,�/���G+�9�P�tZ�&+c��;����Q�T�(��o�d8����^L�0Ȃ�tK�l\��(P,
��n�Qe�A7*F�'�ꉻ��ɀ�ŷF�T���+�(>����f~[c��L��*0/K�[�z���?V�OA��xw	G�Y�Q�=�<����xy��L���̼�Y�j�-��h��:U�+��o���"q�+�k��a��1+���(�	ޟOY6&�܇S�c���b���m�e�>T�;~�u��
���\�u�=�x��߿����>�c
6�ޛUD�ޮ^F2�����#�"�t��;��/��T�?�o�0*�>��T`]֎#V"!�����ߡ̛�M�ko���=��	C&gHX��8ܓ�d#4�A��5��0&?�Z�r�E��i��
\X��_h���8I�����.#.�5Q�8M���?�>(�߬Dq����n��ߋng�s͙o��N�݇�0D�y�v�HU���.��G4��� ���Y�#�TѾ���\�,���Z����Cj�9���Z��y�lMC%e摵c�*�DB��h9�V���@ͤ��C�WQ�$���bt�՟����qT��2����vB���֧\�6�	��.���;�c��$�iN���g�ͬG�5L��O�����e��H@E���D��*�������}$����m�꘎@Uf�j�!��/�f�m �6@����޽JQL�tY��{sL�f��bݛ����&?h�dԝ	V�y9�5�NӋ��~�^��be��[,��5����~�A���S��~�Ĩ3��e�~�v���'�52�����K��ꆳ��|���31T_*���H�̹ʐ.�Z��ڠ��d�z٠r�o��˔O������ Fj���U�$w0��:��Z�בl�*s��` ���=A�T�v�K,�r��#ą!ؽ���p���d�$/r�5�",�t��
���{6�Kv,�JF�!$���}������>�G�c�5�1�Q�bQ�g��qA��-.��� ��!F�ƮX��1~�u��G���2��F�\W~t�"���\J������r}rB���5	���V?��xb�&�#��MخVj�ſ�5�����( UϚCK�_���K�5]&�$Y���:eo�DS:����ip�
�{M���=�&Zm S�n��Ɨ��8@u��q��r�-�6�>��S��_Գ����㮴�'(�e#��<����M8�X��i/{�Q���t�âKc�����j�8۳����[)X�>���O��o=���J���L���r����\�>��!hF��Q;�\�q`?>J��w�ʪt�i�%�;�p�8^I�t��-=�aR��o����<���k�h<5R���x���j�Κx|�?����pm�΀>��5�r�മR�p�|	Y�ү�%�@���by��]t,�ϙU6 ϫ�w����,���@��$�"�q:	m�fFȾ��ZpNf8b<���/�jM�NLÓk�]���.-'/��k����Z�/�@X.:�֍��(K&T3�&�]�Md��啇_�.�.��8y�v�r���7��c"�k ��Q�G!�= ���N0g5v�:^Hqm�E����
�Q����0&�P)x�^'�k~!.�G�M��بN5SA^I�*.�s1�t�;	�=J����R���ȁ���=g΋	_�\��#,v��[�V��[���1�29��$��t��@ϟ ]��.^�(��M���z�<B⌞�$�Z�VqS�xS���JfMhg��Va�F�Aj��G��Wu���;��'��*��^��PRX����sU��.�q\�% �F*�ʾ���Z�x~�K����t���\0d �)�#����d��D��f:] K��R�������$M<����5R��T���L6Kn�_r>�M�u2�Wh���<�%�Rdւ��G���,����xڟ3�o�ҙ����h����m�/Ұ�Z��ǁ3{�q���^*��DsfF��8�C�w�k�7��$��,  � ���j��Ⲙ�y0�W@��l�n��I�f/���~+�X޹�p�v�)��ɰ�/f�1}�yQ�w���jA�#|���:n��]nG*k�l�$�X]FqM����2�[��A�z�>v ��!��߿[�����q����Ȼ��FJff���$tZ3�l���r,1(������0�V�7����qܧ�EJ]�`�o^�P�8D�2��]o����c��S�xI3�֒~�
��+�j�U<eo�L�)��Z*����ƋqJ
$�n�=�8��	���>���R�V���LD;��7�۪��"g�ePHѺ��S�?�f� ����|B���Wȯ2�E�Md����i��F<ƥ�4�J�M���D�@4k�k���t&mD鮞�W)���9<�/��C����O���v �4��v^_'K�%̎t	߾�vWZ����)���qg�|7��b�5��{�ą޻$>��ƛ�K��P%�F����7!��}�6�R����&��Ϟ�U.�(5��	��>��_���"'�*L�>�H����rO�;9�o�A1GV��i2�`�gk����	�+����G�7�oR��yu��*�#��r�� ��v���U��uR9I�N�|�V����&s���}d��"M�L׺����H �V�c8,Mdϋo^_�fz]���WT��M���D�Q��K�J�
�n��D򖯡���t ����������!<z�] 8߃O���G�ڪ����sh\*�5b�Z�ZS@cM�[��f5����Щ� iE�X�3��o��?��?�d^��:H�Z����E;PEt$[������$(%	�������rCn��<�I�m\�����9��Y��D �R����/��YJ�� ����L���K�Ǽ��ċ�.>�%|�*�d�9�&V^g�(�P=5����s���'�����.�W���$H�y�#����7d� 1~�Xr��u8.$���85�(�����3��&w��Ã��`���O��5��G|Y�q ��}b���*%��6�!�E(����c��"J_���Z���x�ǹ'��Ōt(�F�z�w����P�l������pn�NCU��N�v��neXz�ev_���X��PPǖB���������">�8,cnkae_u�9F���i�}�/˸�n}?!�S�{Զ�Ȇ	�������h��c���ў���`���Ucۤ�(�6-K	FCI�3L6��H�}g�m�{���	�O �y��;f?
�ƃh�BT ��~�a�^��R��&�z�_�������"�!��s�V�T� ׶g ~����Xg� y�j`؞@?T���0@#�^֮�_`[!����8駙~�i?���v"�1�[�����%��8��.6=7��r�i��<�hw�&_.0S��:�e@m]���8;>���YE�.[
��p�ǔ�p�㰌���e��o �M������IO���G��N�Ԫ�	n�~o�w�o�}�k��?�������E䗱,�u�e�+�?�^�����Ok��-H�Y�DbY��������6(� �^2y�'�t:�HG�n��� CG�Zٌ>l��5��� Qo��R� +&�4<��;@5P�����e.z��e�G���:?0F_d�m�Z��c �i��V�ד%2�г�䒻0^�:*߅��ͩ�vAw��@uĢu�e�x4�Rֆ�VOY��o�� ���~Ў[���?�F6�x��h,�����0	��+��݄SK���-�[��qW�YĮ`�8�~���Zl^N�>e2��QY�ڢ��M'��3��N��5S2���z����:�x�nq����اp�9��ח�p���N5�E��e�{3�\�g�p���T`��z��tO�M�ƹ_����09�.�WC'�[�aN�y���D���ƀ��0��ѓ��H\u��i�k_uX�q�s�@�tB8A^[��MFW~��"�xt���I7���/�L�ȏ�f��Gj*��/ča)��7���O��A[o������
	���#,�.i}s�,?��� �6�Y�&ՠCٗ�@�C���?-;�����'8lo8Hۢi+���GRg8�=1z��� ��s��f	LR�X,�;�9��,Ȅq�cGo�ɤ>��>�1�6��&$���,<\�*�e�<���F��[�	�da�� ���ʦ��P�4���MA1���u���cڱq�"�~q�Yي�㶄+��\�{̟G�e+��K\�[j8��E�9���{�˖��eH�{���ͥ�fo�3��ib�h���ɤ�{�W>H�Y�6�; �w�kq�K�ź��l�\l�\�S�(��v��H�nbs��6�$�X��\&��	G�j&��;�f]�����wKI�5Z���M�pK=�:z(����ªK��Λ40pί�U Ŀoϳ��z%/=Wz�1��������*�j�"4����M��
ܱ&��u=��
��3����H��$���n�o93>��b���J��翣mc$-9�ퟶ���6�ԿM�+ ��ƞ̖��pO�Fe	��q$�2�`Ӯ��N��ן�v��="��ȾS��[����4��I0�tD�4�lY��A��7[$p/���n�Rw��c2�:��f�E�c2l\�G���J��{�g��u�9�%>����A� . ���U��Ĩ;�Ǎ���վ�lY>�}'I�����&
<��r �%�yA����|�w�NO�f����^W�-��L�Ӭ�?�W�o�?���L����0s�]�M!��-����$V��>���G�C$��IC�h�Fܰ,A"���� @W��_֎?5�(߽�i�Q~'D��q@�=	"2�0��2T���l�q��NL�����4�����i���f���٨U����5-Ŝ^�wJ�h5_�,�B!�o�-��r	����;V�Q�٠!����9���1XY��G���a#ٓ��ȋ
�Oi��b8�/�<�EY�g=����[�)��L)�o�t��U��)�3�1�=jc���ET��B���cn�E�`��?�i�=	Y �ԐE��'01�S=ya�J$d�)�ͼט�G%����c�W�D�!_�ƜH3O"��������h֠sM$c}�k��}��(�!�Q�cc�/ f�/��Uhٺml#]�87i6��ɟ�-]��;�N�zJlv�	f�'�1ze��=�;����P�e�6�~�oh�I:F(��R�CRq��� Z�/�_s�P��1&�]J���Wܠ%��@��[1.��+�=�/��v!���(Ll�|��d��W���1Þ�KȂc��z���G�3��@a�|H�t%��w�b��*'�k�2/Wr����fȐA�[tkTv�/�x����+<<%`F�iC::v<�>�Q��~A&+(��E���03����6�6pA����`b?���9М�W��Uz�T��Ha����y����Ѱ��kB��B1Q����8Mң��&�����Z�'��Ǯm���3
���{�Mk�����t�פy���^�$SCa/h-z�0���m��g�O�@MU�|��?�`��_�$I��̓ד]~5[�5�/��{g�G:s,���r��aL:Y1Pi�b⋏Lٲg�p�p�=���?V:|ɁRo��icҵ'��l���=�5C@�o�t �uT�Fک��e|^]��� B�ቃ��\W��a�Tm4�s�e���ܵ^^�>.�孛.���~>�F��syhxp�9����Dr,P�N��,T
�gR�(u�r�j@!��}��}�&�N�M�g��$^"��`�`�[g�\�����~��-Z���_���W� a߿ʄ�"�s��cY�/�x!V4�8��\-(�>��	��9������J�3�ڶ �ۊl���O?CWVtY��l�(���F��K=��f����@�.����k�ՁEf|n�GZ�ki� =��N��Hv?X)�l�z�+j�C�!)ϸL�d�n�ǳ��/R:74m���C���	����}o�:n0���S���AK�1����
 в��?Hҏ�M�AK��j�v�O��Q�gO 0VA���cv��7�� ��~l�����HOME���M�gM����;l�+�X�:��{�;�x��*o4
�ML-B[Y�@�.����|�;LՃ�h4�<�7���>�=�<�o�Q%��<^�i%�'O�xK�W[%[�9�u�h��*��-Z�T�̧PD�@�d�LQ�ӪS.Kw�ًj��}醉��2���8��9�x�X�~��0I
�р;hm�lcfhH��q�r��b��V~jW������>���bG�Ҧ|�V,D��Q�zfJj!�@�
$.H���&��h���ƍZ�Y�.�	��O6�i�$��5���(D�S��5�<�C����a�N��99p)��뽣�>LfP7�(�^��`�c.I,����4/�i��Z�U��6�6��T�v��<*uW�>�3��^��T�H5�1ر��O�/c�� ��/�f��c��rx�%��덭W� �3iY"a��0\L`a�<ѨT�'�n��.Io��T:���y_���@*C�YQ�OM:������b8�4�$�O�R�7+�z���=j�׉J&t:�+�a?��A����p�p�������j� H��Y`�Dֹ�����@'XrI2�`�C�4@�'��. i�����W���)�jb�}4�uwx��+;4���U���I*�Ǭ��ؾ��^�~<5�>-9�
��T�U�׋Ja�8V|��.Xm�l˘�5 ����o$ľo[�Lƀ�-o�ͤy߷���J]��J>�.��a�)}~e�e��P�dA�c��}� ��Lr�̅T|ɖ]/Y(�C2�h�Lb�rv!ȉ}��>��z!�L��_��%ɑ��ú�����{�/��[:�'A`O�~�=_���'���3�@7u[��V�@���뿜D%��`����=�#8�_�N�a+�j��F=�*�� rjn__,�?��tĺ���#��_���>�M����ht�}�F��hñ��w�Ne�z ��ݿ����^�,����ˎT�����,�k׆��
lu��VEr	�M�qu}:��E�{��"K8Ǳ	4y��i@_A �����^F��R7�AZ*"a�M����u�#V���@d��
[T�.G��g��8�5���L��K��H|9ڍ�'�IX5��L,\���Q)Q^��@��B���,%1r�#�W���k�#]�p0 �^hq����9�ss|)�#�Sſ���RM��PԳ�Z��� ��	^���
�?�����M��vO'&K���S9����J��I����� l��~[��#�B�8	� v�i~7��:�x�	��D�e��xzG��B�B�IA��UО�+rE����ͽ��X���\zy���%#�? x�������23diI=i�L~� A��n�V�ۂA�sm��@���ɑ�fß�ݔ���V��)����T�z���A����qq+��'j��?OS���3���3�&qJQS�CD+��8_���_==�b�b1�/t0/9���f;Na\NG/��;��T�����l9��S{7�틎;*��*[rT�ط��5U�<>�i  %5�D�����u� n���?g�S �ش[�ozb���S�U�%���-TQ����F��}�(!k�=��������5t͇�u�kL杒���+�����F�{?��8���,���M�fr�u-��9����*�"��ȍ�M�3���w�.1�ܿ��MW[L�F�he�;��P��+�������$k��;+&�2(	bꅝN���R�%�;J|j7�ES�8�������<��>Q7J��)�QJ�K$���&��!224�YR(���U�bF���hZb���롶օj�ڴ����
��f?�*Q���M��Ywn��d�{��4}�0��͘/�G)Y�1Oa58���v�oMH}6H���:A� ���F.�wZJG��	aP�VY,|[yM���!����[�Q�h��Tġ�G>��l!�e�)2o#�2:!]Ƴ��Z^�Sy� �A��J�8�kU�s���2��ǯ�N�K�O�E��rUzG��^<�9�/*������O����� �Č��$=�m�Z5Ǝ���+�a����C�#g�ns��1r%J.$�1��>�A櫟gZo� $D�	�I0�
F�i����M��&ϕ
c�i���89s�1O�c]���&�^Sk�ƅ�3x�� �5
YN�ܭAC7Љ�״��dt��hG�6rt�.���7��Tr����V��=�����Y��2f�HwXlxV64EB    378c     a80ޱklKy��L~g(�x���f%:������� ��]%#2�z�!A�^g���A�5�]�������'��>�~ԍo#LQ�Ey	���4�����D��q4�^΃=(yy��FX��`�7��^f+�l�?��o.��!iv0B�t�
��)5�,ژ��4r���Jy�M!��{��Koz[FS����ʎS�]>��
dw�:�����������qf�i���������'�������r|[�(�W?n>���y^�nВ9��9}:2ՠ>��TU3�,2�yFB?j��KM�؉l��O��|"����A�Sѵbep�ʎ2��ڻ.M���g�]��o3���&������<q	�YUO��|Bc���n�@��SD�� $��;�6v��ti@:�%G|EJX��q�M��r�V+)�18 ���ׅ���f@؀�w*�p���C�4w�w�o��Ё�c��1�����x5t�~�1�RZ�����Bu:~X;�P���ꔝ��JM��c��ȇ�S��"��Z��P����O��]|� ����u���i�VȾ�1�	?�ќ�Ǎ:�,�B��Y��H0cE�j|��lI�`UB�F���Y�y�i4n+ &�J���sxfH��������}�C-/x��;��rCz�T2��`x�s3WIG/=a�D���&�?�mL����wHwr�M�N�8�]
:����������;����}��y�Q�3#D@p�Z��CBK#̄��7��P#��?ls��`3=��� �	@����=�7����⁝���ˠ��&^�]�8��l������[���H�Sy�7}h�4ʢ��SMM�^[�t�����T��_��I��Cb޲\fc����J s�!�w(�]��B�I�3TE��e��Oܫa�5#�BV�c�Ey�{)Jh����mu�Ύ��6�\÷�3TK��h���-9��ԡGI\I�8Q��2NpQ{��Td����p񃡮���쎔o�0�'i{�����|�:t� AK�xh��N�d�Uq��G���/ɓ���iK�."w�����JEb�	uqos ���lR��^�L�9�U$2i.-���6@�%q9��&U�ϸ���?����x�Vmw�2d��M�ഡb�2�0$p2w�c��,V���������-�H��$Gz�2�5u�>�u��eǬ�����^�ǌz�����k靜:��� 2����-��A�Vmi���07�I�=N�v��e��o?/�g����2�f� �Y{E/W�it�_����/d>�&���
�3�F���w��{쓤�65������LᓎvX���__%��Td�Q|���� W�X��R[Q������3C�\]"��0jq�v��"N�����3�iT���(<8ӻ[��j�dK"v�:?�D-Lҫ'd|�M���J��b����PZ�jf3�7KнE��&ӓܫ'y8���!A:�ϜH@t�mՒ-yS0�OsA\��&�h�a�M��_qL����<1A0T��tӯrNM����aX�U�}�4�a���A'=�5d�s��~��ݤ�!�fV��7裝���n\�o�NL��E�8�l�|p��M�Z��QB%����ɓ��J���쫟�5�:[$g3�ݒQ�	`���L/qɺ%��_��4c?�ּ���)�����?zH�����Q�]%�XÓN�H�z@���_��-�~����W�TZ�"@�.�޷W[N����Y}���hؒ�朕~�*6�|m�}�f���RT�:l��`Q'1�"����Ё�q񰏖�8En<�������"�����ɫߥ=�M�]��ӘA���ނ�t6�]��c�,�c�q
���C��^Vg;��С�+��_�Z����kԭG������ӌR�2���S�J?�v6�/��\�ΰ��r�d�u���y4�^�2��c/�{�[[/~ox��(W~���""����]7�2�jM�&h��[M��X�t�v͖��S(8��y!��n�;{d��69�8[ ��F�]�=��p�u�J)I�v�]�]3��l%|B��?NPe0_#�
�TB����3����1��O�����v�7X��*)��j*��X�S1<d��.���T���D�m��bp�
tn|k`��:��b��m�Z��	K͛��Z� �вWCx�ˎ
�Uԥ�?��-`��i�;>�!,օS���+� ��C��c+}'�4=�[�!�����]פ�Y�����s��Ĉc]#�*�P�ar�
ٛ�w4^������������U�G}g�%p��	�ӽg�7].� ��:ϵQ��)ՐZ�d�Ǒ�p�j�X�	���I׍!��b��� � Lr���AK�E�	�ള���urL�8��a�U��䳚���I�Km�j�9�n�n���Vl|t�j/I,���,�|gJ�P���u��%�Y��
1%	��U��;�\��$d-�nZ'���1�w�v�֊@�(����i(��ӕ�"�'�*)p̠�����V�C�s�d-�]a����y��nuP���d� ��/�\k��Nxʳ�)�T ��a���
�$���QÏE*9�E�Ƙ��g�'~=��$:fO�>�����kLZ��n_ǽ�"c��`#����