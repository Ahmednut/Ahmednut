XlxV64EB    2d58     a80����Aݿ���ڧ`��lV�[�+��ʼ����Wh
��B4�,m��|���!�>`e���b.��hEu�e0��x���$L�D�o���W�%cǈ|70t�%n>�ִ
W����ml݄=+������wʶYM����o�%��< ��ظ��B�{�$"|V.�fbȢ�\�Z�]Q@	G�߀��<�|#?u�0��֜�� 2JyK�&�Jk.��Z����~F>q�������b��".d8P�h ����#ۈi����h�d��n���:O�a��>�2�ä��Z6>�!�噩����w���C�A9:�Z4��h��� �1]0�p_�}��J�T�Rp��P�Y��%����a(�gO���}R\��i���l�V�^�
h��SFlE.e-pvw�?�?P2���~%x|~���c��	D��\υ$���J��:U.LmD����muM$ǝŠ�Ҥ�U�3y���($�H2��*�ϱ��(C�6��o�=��5�����>�k�ukW3�T�*��f�tI����G��蚘ǁyjt�ʹI|1���f7��\�ߖM"�Ooz�k��8�����,S�f�vx��"�k,?Hؑ�!Q��7�� ���a���F΅`9�����$�찄2	|�m]z�`��1�Q]D��7��wT*��U�d]a��yž����! ��*�Ru*���������Y�Z=����6���kj|B(�-��Z�O3H'da=+�Fx0��jԨ�3�ɔjg�a�������ce�"b`�I��`�*����f�6�9��o�:xM�X��O�|�&�[����F���Mk�}� ��9UR��d[��=������DRP��1��o34/v
�ii�9l1�ܳ���)����9�%I�G�Z����6	����u46Ʋ�'���o�x�.����y��o�T:����R7nc����LP}ϓ�x���l�	i�&����pkɢ�Ղ�z�r�I�jY�G��e�N� ����Y��B_'p]����7��z2�gh�\B/�W��W>"/1���`#j��
Bk��u��J\҅�@!~yC���)q�8M	��?����Pkr�ή�26Ic�d)e��g{\�h��[F��)��\���� �L�x��"T�����F	Q4�������0$ߨ��#�H��Ӭ=�p���F��K�������WI�a��I����W]V���[U���ǃL0��A��R�p8����d��м�ʡ{�Y�uW�BV_8���G��-�:h��WA�NM��h��ȡ~�蟅�fҾ3�3�Em���4e��hsډ�`OX��|�T]��Z+Q�>��l���`�غ�(�&�0=<�z(��v6Wʰ�-�7w�"/�a�u+��4�Y��i�F���+���N�L/&�]{�xd��H��]��p�M�5MMM&d|���S�qô��<a�$O�l���	$��Q�A�� f�rk��uP�\h���,�f�%��o�\p�OJ<�H=\��.n�ֱ�}z&L��Uj�1����4Vжƺ�Gk�E&���{x/���9�������3���f:� A���,1��U��H��LP-+�X�]��Cڂ5�����Wp�K�)X��|3�=&�^��$ך�<9�)y��f���?uÆ������N*��i��i�Ft����,�6�ƽ998��t�����8�,<-Y�2}}�WL;���"րq�g�n�l��a}�%�*(`޸��z��F�� Ś��I��3��oH0�O2�f�axX!���ĸ�̽	�l\�-�I�c�\z10��i):�An�f�s�Я�˨�E{���FQv��'�r����(�Y?V��|�ܟ��M�d�o�|�d�f%AAh
b�,pai0��B��[����8D�Λ�v�m�^=DR�)D��?���$�n�o���)��q�k M+���4�ؐ����*�n�w�:���Z�}�N.\�a*�Y>@�q�kAc��xEt��0`�նU9Ρ]@-Dx���0�S��3����r���!�(����}�͕�-�S�]����_ZJ���:�Y�,L����g���
�[���-��T��Ւ{�}����p����_&��׌�rp햇-��c�'����IcCk����
X�Km:�/��77m�]��G|$T�%���EK7����s�7�eh��&��J���i2���8�����8�U���>	��{�#�E��
�H��Ǹ���[4�
��}l2iS �.q!v���	��?kV�����&塶E{�G:i3�h~����I�Mjw|+�#cFrP�&����tҍ��a�M��?�!�dT��C�E���ML�D�,�}���a���ǿ�	%A����Z��1�Є�8e׀Bڵ-�>�zҴ!3l��L�bO?��d���>�%Qh[p�$O��Bw��Ҏی�+�D�|����@4��;l�X��Xg8��8�؜p���H�m��
�}�
4n[�ήD��_9��S��o�����N}��0��P{��P��G�|#�Lg{Y�k;S�ސ#���pm���Q�/ր�֚� ~�c���L:ߤ7Ȉ�`���!Q�9O\H,3ČZ'�7������z�N�P剷!������.�T������