XlxV64EB    163e     870�
��w!O�sP_x���y<����ŵ���Ij���wn6��8����b�F�N�\ĳ��Q#���=�&Beϟg)�mY/ζǴ��(Q7���4Sq��>}X-�5{�z�H���Z�#|}$n��S[��w�����48���	��Xke��(���r�]���$n�*�B���0]�Z�5�N���TsPn���9��m�[�g���n�s4䍝$ּ8A�b��uLP-We,�	�?�Z�;Bďz�n����!Պ���_t��w��7�G�8l����qٛqM��J���ڹ%�lXc��������>�	�A��8��6��I�$���s�ɭ�S޾R�%��A�dDL6�w*�vt�`&Km��g�ᬦ���lNc�U!�'����B0��$���]���m�q�흏G���t*֛j�4z�P�'����H;`M�y����%���9aϏE�yO���v�?ɿ~�Lv`�<>(���i����D
� �b��i�ܛ�7&,�o+���u����M� �@ �����R���q������+�>٘� ���,���MD��ZqQ�O��k��r=
��[�E��  �����<<��dhy�d���]�_�P��� ?���		 O�8��)Sjԣ���댢Fa����z�T�N��v��$�q�r�rZ5`�R;�w+�B<�=G�n��ݩ������_���)%���]ϑ��{��®��$��ڰG���<V��+���$�'{Ƭ�'�f����
}��S��(�u�F�;�A��CpETy ��<Ј���<Ԍ���=�/��JQ#�8I�h�e>[�V�/�-�猺p���q�wy,���a*�:%	�[���9���P>�E�H�_UfF.-����\(�6f$F����V!��qߙ
�l7:Z`h���E��~�$���/K�����x��9B��(��{����E�k7���1d��X{��t�L�Ȕop1�ʻ'隩;F��
�>��.d���M������-r��Ck��mf���,OGx�˺�N� Vi��=L�!�Y�i��>=�s1�mp��4����nI�	����{�U�����:����#���^%J�r�=��G�v<o�u��AX�EQ(�����7o����o�k��Wk�pd-�_�N�Q]��#��7��� B��}���Д�����~�?��naո>��|Py�p%Æ�����:K��[8O@H�;�����6ׂ$ &
���j�c�Vxs���4�X9�vi��׳B������������1?C�\��^1�G���wI��s��`$:��Ұ�������(([��Z\�Xθ�z{�gn����4����'��M�ʐ��-!l���A��)��e!�ː�^k1hGl�bq�L�f�#ˉ�hmJ�^�
$g	Ч�D�^M���#2����Ӡg)I)��3��	�5�9��FG� jȮ�h�`{o���8�&�O�A���Dq�2�Ɵy�E�@�gx����g��b�@�����+'�:dt��"ӡ������b:Zo�L�w�Kzd���B���ï̹ D֧�k}�0����f����TW^��rk�2��FqCM}�1��gr��˄��~��>yXQ���~��͕��"�V��0j���-GW���f�"(�kR.m�W�g�����0b��DLZ?q7_���-�0r��$�J�7���:�Nq�Hv�Y\ft���:��}�[glS{�s�"o2�0���O?e}mo�� T[�+�e������n�[�-�0(_N�~�]�_S�ai&�����p2d�./P� ��B=�"�M�v�UI�~B"3�|
�Zk�
��z��"�\QO��#�����m�AG
v��Zړ���tW(O���m��#�aA�.����SH���D�����yS��ט)��E��$u�P�TH=�g,�B��]\��b��I�9��$�8L��1��Dl,�ME��HU�7?��K��ݦ�u���Nũ%&��l�½3@�o(g���A�%VHA��1�iՂ�]��J��Y�?)�R/�ц=�i�фV�	
]�c��o8<L��%��{3�l��}\��i�:}S-vS�������O��g��ĵ(����m�*β?����{