XlxV64EB    1945     9c0%����~�n�D�*��\V� &	��W�y;F�f-S��[w�+�\�~tpЏ��d�h���a�x�}��=��/�D��S�cZ�
�w��d��c�/��9((@���Nf�"��+\�e
ɘ!Z{����i�)�8v���iRdc�����N�C�4ʻ�e"i�_�ĳ�(��%�ӄ���hŠ��JA������΂X�TBK�+���I��g-�Dsܬ[A�&�ꫨ���)�{��,Ƣ�:�>��Q�����٩�1���X��gŞ�v�M�"�^9թj?Ǣ�%���?`9q�+��]�W�O]2�2�3�׬��#-�-u~�p�y6"����
V	+E�N�*=�O�������y��JN�.j���^����G��K����n���@s�E��u�bח:�ݿ��L��x8��ؘL�-�by:�&��ƛTpJ%o�0_4������M�r����v�`�a�^^�H��i�ʼj)�m/�M�W0�*����cR�o�Hy��w��ٶa|3u�瘨6���E��@y��ו�L�y:��T"$f���}�g7��q���xawm�m�劓�� 0&�Tќ��j�߅�y3�ك���S��DV+")eͻ�7�W������vYܶ�n�S?��|Qg��z��=~�.�\��'�ڡ�jIJ+�O6���G����<ʌ��d�
��5���<�5� tƮ�t��b���£\�n_�&3V첞�5�3ד�F����x���8���N�4�_K �2��ô.�YI����)�bQ��4��r�#楕��Y�;H�����k�%�l�O�	S���{�~�,9"�t[Oth���Zw���Ӥ��� M���3Ir.��n����ʆJ�T�*�h��my��ФgLo��[�h�ʙ	ȵ!��n��B�Ϊ����HV���?�톀�Ż�
�&�	I��AKq[�c����L�'����0��JQo��Ϻ�&��qF=�r�z��E��|�	��!��f�������x2�l=mt�"ol��D7���G�t����Y2C>Vg�p�e��[� e��c�n�Ρ�c�-8�eɏ4 !�p&c���e�7e;��y�G����r�8�JO��5z��}g���C��p��G�Ŗ�X�z���ዷ�kOc��>��ʠ��hC[�]�)�RFhm�@���
��'��ІV�k`R���m�=�),��载]e�Q��Tt�W���ōs�T���=/�6%P�Uc^�D+;t��uH��&��c+� k��8(v���HV.��o7�;�����t�	H:��*N�o�_+��\���1_����vO�Rr���Υ<��ŝ�t�7�IOT���W���>[�T�&ѿ� ��X�|�uG�-��]�٘̽}��=ފ7�Vj���7*�g�������NsTV*�/�
��i?)���Q9�;}eܔzT��f��U}i�W:u*5�c��.�9K�Eq�(�K6/�jk��	��h
�[�*ǐ7x��u�v���������xAm=����.7��d�2��	�XF�)�5�G ^�Br�7�S���g�Q��:e��}�Hq�^�1�0��Ə�t��ۜ�܎���O���G����/���{�*��X��vP��)��p��+#�7���<�h�Y0�?<���t�C�G{-<�d_����k�Ip�s�\��-����h��^e�o��IU3"ϕ0�$�jJ�h�
25Κ��~���o:���$���P�CT��C�:�T�Pd�
,���������PFx�D��Ϲ�9��:}� ����U��@��_h~]L%��?6��`�j���K���,��|�#���n�����~ə2
ٕ]C��jb�����Ά��q������ø��NLq^<F?��B���
)�J �βW0��C�%�ݲ�F^�q�"�=��������1VP*1�n_$�G���@�b'MI7$���j��M��L/�?��D]x�)�����L��L�.��� �,�e��S�%�Q�I��H�{�Z���zά�����a�8�F�vaNwfm��ȗ�ᐉ#ҩ�i��q}�lԇ���/Ђ
�8����|�ݾ9]�� /���oΫi&���"��/�r����t�1�?�X�~d(�����<X(y�����l | ���t4
;Y�;~e}����'xZg���~Naʪ����<�RS��J����C:�P�p􍏧_0��q�L�aD]�t_f��|�a5�Q��j���Kp��+՚q����#v���T��b���6�>�S�ğ��%h�,N(���V�d��Ϭ�hL�β�	����A�W�G,Eg� ݹC��prv�+����� @���;~��lْ���Ǽ�%�Hܐl*s��U��ҫf��,쐓��]c`�u�<��0o�~�c�{e٨�EU �G