XlxV64EB    17dd     9a0L����+m1��k[l�T �m��=�"��C$���ӆ4|�UZN3��QJh����z5̈k��{�^�F��Ԓ쮥�;l|(y9ʉ��;���az���9�;zx����1�����v>w�g�m7��˯q�u�4n\N>�^ak�����Ĩ�5�?4��z�"ئ�y�ư<l�P:��T���$�g3��:N��b�2�v6����7O,C�;󣃇ͪ�.gv����ق��of��H���\o�+K�i��8v��v���r�(���~�d��t�*(gPs�����cr�6Ǒ��� )z�_?�_f5r����%��I%��I�
�A0\)T�$;$����_���ڭ����E�h�I�}}=J����y!`p��Z�i��N-����ʽ:WVԼ+z�Xk?�f1��U����n1w�o���]�q�羲\W"!d��/��l�����ƚ�qH��bH�)^�=E%}̏��L>��yzR{D��r�&<�	�7�1�YLL�1�����X�
�Z�Q����,~�2���Q ����0�?�LwR��K�ܠ�0��|8�EHo5l\?=C�j�r�/���i�0SL�*MB̴���>�1<|��!B��G�fyWY����OM�8ZId�a��m�nr6���#���Ɇs����j`��V���]��9ʔ)�)wvb�!��8
�dc�*��q�sw�i�@���:W����.��L+~
kt�!˧S(5l6|��X���.&�G��[.��@ߚp�����e���cO�f�z��-?���D}ʊ+���7��R����kl^=2�K�8���$�2!��?�F�d�8��~M�4��!��%y��.�02m)(O�##��G�
J�cn��sTۀ�wx�M��n1�?u��L]l�.\dk����T8��6��e���_�\ն|z�H��"��\r�^Yd.E�|Y���Ve��RxB��Q��Q�a,�~�
�1 ���[���o�7��,>YkTP��D�$[������k|�����I�P�wk�EKQ�nH�� "cr�U�Xh�q!�	�N��G�����1P* f�n������j��^3"��8Xm�Rj�T���c�H�2������? E�}D�����S{�b�V8����W��<tH_x9%�@�KR1��'j��ZW-E�)J��5x�[(D�P���B��@��v���RH�/|�cDF*��eO��Yy��Y��n�-Oe�1>��4٬����N�������F��Kؗ��6�g����)�%ݸD����XcCR�`$2^�%��vؠ�����e�H�H4�x:�1�! ���{0�"4#�����	N�U fZ}�L�&�;d���s�֭I���#��Ŏ�,��������(C$�����6F�1L%�2=�6.�Y����Ü�6�li����(�k:[�DN�#��T���e�X�}z��������@	֡y~���f� ��/�a�2���|�9J��iȊ)�.롂��/|�>�`4^����aܸLL�МM�AWɌ}��m��^?4.��;/��D�b��eVc��z��3[���� EG���)��t�g�\n�����hӄ��}ᖹ���ҴD��T�Q�4BH���Mc��~��k�;"v<(F�kZ����� }Z�BIB�����GC��p9P�������j�Ĕ����\�%�x�1US��(_��.4� �#�s3K#"��`���;֐�<�F�xy�w!�9+I'ھ�z,������O�P��)���bw�(��h���*��0`�)�]���.X�X�N�>i�k�C��]�qB0W�h���q�
Gs�[�0r��1J*��a�ф�?o"Y�8�z�Yak����pC�|?+V�5S.%��P17�7{�^�D��h�i��dipG^�(yE�_�h�<�Q���z4��+����d����ͅ�4��c�~����M�c�!���B�w* �(��!����)n��&�\�X��!�]�4�;y��!���.4�s���X���ot��L�������"?P7��
w����t��EԾģ��>�\8��!���c�S��@I��Ig�w�^�..��$��
��9��e���\�ӑ4�I� �r��i����l�H^�t8��& I���3��˳;뇄�pߨt�FT�:�;y	�j\����B�S_b�|�� R��4��=N��#�߼toӕ"�b)A
I#w��Hf����f$GT����k��Z��:.1~��.қ�ڡt[5a��Kv (��.�&������8��W���
�m���l��U��v��?��&�M�X8A���ID�Q�Z�Y0e��:��j�>fZ�����;�{��&�6d��S[��<��KWI<!{e4tJ�&/�O�