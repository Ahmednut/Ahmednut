XlxV64EB    490b    1160�5���=�N���Sؖ�����è�=�[�ڸ��!�Hb��J�h_`k��7r�+Dz�~*�c �v1��W���d؄9� XH��� �m㾐S[T�H�����(k�1��õ WqN��A��N��g��0SqBI����$����a!�n?�cSh��3�*z%���꿣J��Pe�Y+���6�s��7��/⤍�ĳd�a
��i�Ջ<.�`���ֻ@d�QI��#��K=HK�ИX O��zk�[�  yc���6� c�Ao��%9wzA.�h�7��{'C���j��arA��}�j q�*�b<5{���������ً"K�������Ÿ9��EU6��S巶�d��KR٣{fP/r��*Y�f�ˈ6`�E��������hH���3PW�\wo��-s(N�
�~���G��yP��e ��׭���J��� &�\tL��0���ˆ&�Ȩ�5���X���2�������jQo�"�-a�4M1\�'�/Z�=M�6\Ƒ�tKS	���L�W jI.���U���p�a��f��R����u��HA�q����	8�L�4p�d|��|�v���~W��Ml1����@U�
�?�����ঈ|�L��cc�)ⶑ��H�n��y}�V�y۩��Y�[O�yϖ�f�W۝��ςmJe���3��K�H�+9��B�@ץ0WI��J�DZ��g92�P��K?� �]�=2�{N�]��T&�֪S��(U6��ϧUup��/�"�_�5-��q�0U�Y� AB��AA�2BGy���e�QW����:E3�䙇W�ib\.F�K����@���R�)��l�/H�1D�x)� ����7aq�8zG���G ��� 2�#����A	`���B¦[��k��sCv�J�Ű����OJ����Emo�{U���u���.y�K�����c��J��\P^K�g������|�+d B�ny�S��2=�<,���^�W�j�Կ>��#
z6}_����':�;����([����f@�tЕ��L$��TD�I����`/�qP�Օ�b�Ig�i;�����5��	��D�h��L�����֙�)�=^����	B�~�����.Mo�|%C��/2kT�E�V1;��E��i��c� l3k3iX��%/�mZ���Px	�x���P�����U�=�ށ �|v�*[\�a�o��-�Ĝ�Ӯ�ϴ��_�$QV�FU�[��iq�ar����+�זo��q�(�ŭ%��ـ'��Ҭ���:?_V\"��8>rbX���F&��^�����rl��ՀD\���\rt·��� ��L���.]�[�v
�~��d���zd!���	������"�!������nk� �2�^�<)��ol�BXG��4��e��UZ��L�[ì��/$����Wa�Q�5�%{��'$*TL<��ʄ�
����bG�� ��6��J�a'�#���{w�xh�2���/��ſ:q���+�j�Z�U�7����o��u�g|��G����v�:5����OO?}��\u���O��}���bՓ�_��6��bC����6�p�
rz�qtQ	v�nC5�@���+��x�#,��A��)��>�$��د�/�_2�(?�0�(j��O�4<L;�t�HʓRI�$~ t��>�:'>�7�L��Ǒi
ǟ�4�CBf����S}�vAP��3���&G����7���>���<���W�`�h̴�^�V&K�,���I�Y�� 0k2JC�������r��[+A|�j��,��-��q�g�ݡ �#����^]cl��J��P;�m�e����k�Y���{ȸ�k��DW��H��#ȥ��3�4��-�����B��>.-��-�0ХDJJ��d
�é����#���?�񨷑V���	�)ਗ਼�A�{]޴z��]���R9�E1"\�� �lb퀈C��D'�r��e�%.��@ES�&e��;�T�_'�Q���>�i[y֛z��@N�(��tH=��?�,5B��?�f|�0,|T玗�9Y�3��k�����׉�v�d �$�GA[l ������#��oR�>'m�J��ĕi���C=��s�L������O@����_ԑ��%ॴ�$�Z��JL;��:6�_t̝iғ~�=̢���A��e)��@���x��VV���f(Z�o������O�I��4���R����Ty�)��uK��Yj���=s��r5-�4���KQIRXa{�(���B�Uժ��̓у)��P�żo�Әl�O�܆����"��ui����[�~X����&����sn(�= �Z�� ��V) �w�� �W,eA
͵�3k�蝭ih�[�˜y���wW���J��y�e
��{˕a�G,��k: h��O�G4Qd�ƥ�@h��PM���x��;�Zwd�b�!�7����@x��U/�gjyG�SM;\$%�4;I�Ψ��M�%�"7����D�JabV�ּB�.^Е-hF��V6�u�cN����e֚����ߵ6s|�Z���p�8�|�Џ,��4n]Waޣ��^D�NA���{�i������'>�T6R��m����p#CK�����m٘߶k��1���x�cZ��ZB|����c�˘��	�2M�m�u�0�����<��k�36���L��{��s� �诎n��7�D�{wFĦf�K�=��	�sET��֠��)��_0�#����Su������{�	�h�%����������q���D��	I���N�CGX����W`�}�>(dҦ�mx�����3b���`2 ɸx����w�,Ƙ6G� ��©0���dw��AM�U�>f�}
��Bfxx_�M�Ѷ: WH���QpI{�7��'�0���RP�GI�O����~���^Z"`�Gn�%�!����1`̜r��ɳ}��-D��� l�%`/��}�Q"�Gu*A���{����f�ʛ�YѨ֧'dv�"�>t��~n?p,�oM���q`%�?V����G7bG?"���hfgY鹒������N[O�Z�@�ge�(�>+{S�u�b�YQ������)��@���M�>m��UO���$�R��swK^�:m�[��,YcO�c�ϗ�M*y�X����F�*�e�©���?�n盲Bk�0btm�<3�p5J�tƁ�f�3�M�*��W~NV=Q�Iz����r�ؔG���[tv�z�p��G8�*l�$�2A_#lD�6�����<��u�%\�x�hM��`z�� $�W�G�b�wz���%kb�<i{�*�'k�:K�G����<�����B�(�6x�Qb� ;�~�YF=�s19��U_�fA���1�oXuK `.;�DSX&a`�3��!��I�_ʿ�.���:��.�W��8b�U����S�~�U~���\>��>��%?�.ٴ�3�=�5�I�ӵ�ޛt�a@L�f\B���R�qxr�Mw�S,�k�d��Y��C^s�Tt���~^X��"b8�W2�/앿�coR��;�g�[\�%�ǵU@���,�h�ŕ갖щi��Q�+R��VQ%�إ�-K�/10 �� �6�*D���^}Ez����j$X2�p!��AR����v���y���c�/��3�~UT]��H�%�WU��\��[�8���{���K�jp?���u�	���,[�TļS=Y~�?������Nc�_O�0��g��� t�������5��u9Έ�7��R�7���u@1m���:NG|�[v�rW>��3P%f"@�������ff��	JX��^D�^!lZR>�
=R +��y"���kN�@}��_�6*���U�������Q��7H�U
��1^.�[�~p�[N������Ȳ\y6~�3�%�Ì��ru����
s��Y�(>=�҈�wp�M��eT��t�M�]��(ۖ��Ņ��ӎ��ɲ��L�5_j�H72ajW�~�<�~d:2��b2�=�;3�0����q��V��^+�ǧO'u)DYI
�\�X��4Ǡ�up!�����*l��M�sD����'\De�<(U �t�|�Vk�>p�c�ū��9���x���<�yP�5A�/��^SSvZf�t�/b�m��z%���ߢ�\�0D������ ,������7b�Ax��_9;�L���PY�~���ʪ��2��Fcj	2��A�軏�Ši*�s9����5�kc�b�(i�Q��G19F��R����g!qx��u��c%߰�0���R�+4��9��8�y\L��k
�}�����]'��٫�qOBW4}g���%|��=�w��W,/']�GZ��� �:Fl�����K'����Z`��E����[�Z���[`祉�CȌ��$�v�����Z޽H����9x7������