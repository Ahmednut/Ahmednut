XlxV64EB    c9ef    1a50�����!N�9�*4}$��cE�T�k7>�݅�9�	t$
�؀8�mn4-�2mR��I���x�sR�b1����VRՎ�ϥ��7�Ag �'B0`^��`�A)[X�haF;L��5�=���7�[��ɛ��������U��O�s�znrX���r����\WX�hsg����܋8B�.p�_�[x�����:l�>�Ú����"�Y���ƀ>����hĮ�1W��]��(���vt,V���ݐ�@�@'��X��Y�h'�T�\=����Ձ�`�c�>qpF���r>,*��t�ǧ�
e�h�등'��T�Y}��m�I�rX���C�����z
����K��K�
��4���4��줟
LQ�1���E�=�6��gvW��ա9��  N��(���PZ] ���w 9���v1���P߻6¦�a�z�W�v�!l!eD�r_�Xl���?�X��f���x�x˨�$H���S�z����iM�N |=6�2�;$����9IM�5��A�&]X���q���-#-U4�of�Q���4�t��2���g��o��{W�v�z�PٱfƳ�`h�6c1d���S���p��R�yX� �.{�2�&�$, �O/�?��g��'��S�7g��X.m��j-�_�6Q�%fy��o�~Q�42��F�h)���<#�+���E��z@�2�
���`���nϴ��|�.��Ȑ\HE������9,yJ��V�e`L��X��5����TwN����ek�����DU��.�ȌM�{��#ʮ����υL �"Ud*����<�'r�_�-ԭ4y�޸-xn��n�y�wNxᦦ�tۥ��T/5��n�L	�:�>w����{�2������W
c�{n�%T&���c3vl\G���a�oV�%W�'�kr��C���%>k��Z����D�%���bV�;g}����>�O2cq`����1��!���1�E|�xm	$�I�	Vo�S��Kx<J���ӟA�^c�s�-1{���p���X��y���)\�{�-V3 ��y �e�%�g��)4�%�����l�̩;����LD��c��\,l�>6r�uA��Y�\_����'^���X���?�u�����%��j�#���A7���y�?FH=���?��u��O��L���P�d6�{���l�)Fk��\���FzF���8_;��Rĭ/��uYrZ�X:���O���8��7/��k�}�c����(�F�s?�B?�r�@4���ֈ�C#�Y���Y}i��᪲DE}�q��3(Հ�3���p�����|��,x�?�[
��v�U�hڈ9D���1�U�z�V����kp{MY)+IpՍd�1~/q���8à����gs`!W�M ¶9���H���D�ʚ/��5�M���V�6Y���|��M�g�ֻ��"��~E�H�g;�
�p��}l���Y+��d�ʭ�Q�g?_�9o�g���,q(֢�;����U����1I�Y�?�$��/���Â�g���kZ�������o�w��^o�D�8\��t�@�>9O[�P�Y�2R�������ER�-�����֑FK��M�"��<F���j��R���X3-��ʬ�u�#g��A��%(�X��
��:�}jhpOnK�c1��50�I��%�?��1-)�vοʘ�m�A�0ަ��n������INC��U���@C5�Ѓ9�Q��"l3����)(��`��2gN�,��hEj�Kp�!j�
�/K*�����d�f{������ˡ1��}�Qb�cm�"���Mt�H�V^��Nq��{UX����dM��;� ��t4�����I�󢮫��V4G?0��P�>�\���6 R��l�-U�x�����R�=3f�A1J#ċt���Uc�s�2L�n�}gˉ��G����.��9�yo�Q�Po���'��V�&8���������0Ԏ��d"ˢ
%�?=�M
0/��3)+�ERv!3���:��^��EC����yP���y����fX��;���)3~�4|aJ�٧��`���������ͣ��$�m��hr�DR%���wRw���]��8��"(��OSөa/K���e�i�m��T6r�q*�a�C� �6���v��B�)��< �H!�c��aa�-#
�4-N��z�~�y��3��ӟ;݈��)����'a�W\V;�m�5Aɛ|8w��D�G�4	E4[�{{��}]��c�S��=l��(��5�⋞�))�� MD���E/�G��h�������u͟����$JH�^���Y�fY��:������,ů��y����(���%,p#�Hb��k��B�3�zz-�X���C������>Z>�"H���3��η��F]�Kd����#d��=��W�z+������!���v���H{P�l~�Ws:8������rQ@��f�ʞ����J"���t�������fz��5g��f����L�8�jK���b
�$�s皛-sf��Q2�µ;E� *_d��?h[O7����"T��wbŔ|��;X$p�}�du�E^���Co�/a���Ul쐾�7}���*�I/�L_<��0"���Uh��R!Γ%����b8�8�6U�`j����롔K�4�	K���]��Cӎ'��������jLX�3_6
�*ܤJ�<����8����3Q��&���($_�c�"�c���@x#��y�y'=&TN���XM~!V�8�7!�x�KZ�Dt[F[���*���˯���������]KM���S|ɮ�LL��pV����u_�e&�
~B%q�d_��L4��.��78�w���a�W���m�	�����/H�g�̈�({������VM(R���{�O��IK�+�=6j���-��;�m�O�����A���S���֮9�Р��R��V:��'/5cn')Y@-���|����lN�&̠����?��,(�>�f�Y��Γ�K��e��ln�W�eM!`n�S�"frI¿��׭��F�������Y�)x�/ۧ<���*�ru�?�v�G�⁼�7{�/ǉ�E�c">��{�i��|�8s�9E8�l���f0s���TT<�I�ׂ��%�=~�#P���1��͑��7�!�WK��._�d�1�����T�pZ!WC���dX�� ���.IɄ2/N��~##L7Kv�v���Y%q�o�E�WQ��%����$ɞJ�ԑ�$s;5�wG{��ơ�(��(�*���2�Ϟ�+��H��W����(X�RB)�Ͽ� �[��f�K��)-�]jj�b��{�Գ*y /���*�Έ�\|6~��Q���7�	l��z=5�]6 !��	?�i��XN`�� ^w����vY�j*�Nڧ�0�z����:C��bګ��Dº�k�9�I���cJ�9�a����Ɍsp��$���$�u���W�P�>C#��	�M�&��������zp"Z5�ا�ol��8[�
q������K���w�@�>�L���(�
񬎧�0���)��}���%�3%�����Ox�f����KPw֩�2��ʝ<�J!v�^��"P������g����p����*i^\� ���`:*�����֐�9�0u.��������(8�Cyr��g�}���
*�Z�L5)�[z���P��|�d����Y�Y����滹Vu�*��-<E���3��v���Dˬ[���Vq��kI��s�N�J�'��-ݵ�V�ÓQ���Kc�ͨ�vD���G�>�t�
�b��"1�-$7�SeIxG~
t>xC�f�jrd�:��"�0�Ni�e�]�^-L*�aǆ�׉i�*�]o���/�z���(ϔ`�7���("�d��d��M�q�F-�l��^��C���N�V Ǻ�C���hq�NpR�$�`�%x��8r|���.b?_�\�ٴ��MD��y�X(T�~0��h,�d̨rg�G~T=�5���ra�3mD��������JK]�hcy��(���1��{"�����xm���6�2���������(d�c$U���*8ߢ(d����:��-��-FTKk.�!l5��Mm@'��4;��y�����E�%Rt���̝/{r�G�Oe�C�X�i�h{�����l������d�z��j�\W�L$R� {�uExy\c����1��0h,�I�=u��̸'�x#���]Hi7�^���L�p,n9���˄���V�s���ԝ�e_�S1�ׇ˕�0���qږuݫLfq>g����a�ߕ�jY̍DJh.�F�^��nn_z�'X��{�x[��:�*K�E�tWܐ9���#C0-m�Ye*��X��Z�3�;Ƞ���0w��<X���r�����go���8qT�7�-\Q�Y�觸�!TAu�bR0�
o8Ah���'��%��W�*O&����5���,+ܨ8.�.����˾7�.'��I�֭��|o+��$�z��$[�!!N�v䦣�!W��!7����e5��'?-5S�8������I�� �R���G؉���&:v~Q_���DLM�z9XO%�4|�ѹUҀ>��c^)��)�X
O���p��wh��27�#�>�G��Ҏ��Cyj�E��IYz�����ֶ*�*��^�,���W�"O� Wh�tu����Z�p;�{+�i�Ğ9_��x7��oz��`��V���� �
o;#F2�}��th,��o�/7c�����~~\��Z ����e��F�t�:2O~���3oBG�O8��?m|�0-�iâ�3�5�t+�������(LdF���Ro�y���]?�O*a�lf7��KUe�7�������m��&��F��� s�<�I�9��S�Xh�t'=S*��� D�����!�<�ވ˦�l*N�g.ҏ�� ��u�o��2��/����hT�W��X/aY��#�Y�5������o�	��bۀUm��ON�3t|FWr�1լ9�l�����e��``�c�V�T��(/�R}sn=|Qm}� ����i�K=4֑mř`J������_��Џ2�	����(��/��	i�J���5��e��C��X����29ElB�-�`�,���sg
Tj��(�t����4�{��m�����x��E�YRh�_Ai�m|��ZAE���N��lDe%�rȱU�m�>	���v+O����Y�X�U<aҿK>K)�s����9{��(�]�f~A�@�����g���篩Q�">F����Δ�q�!Y Deb��Ժ�IS��JW�'Њ<�3t�ui����	骰����d�Y0���Hwn�v��3�
}x�+*��@x�}pA:��(i2�*�rc��?b��M�y�]�<�Y�OiL3@�Eh���0F�w]��,h�w�:>��	�'���+�&���mX���B&I,&�t����v��ca�8��d ��jc lƏ"'?�
]�]J��0�����l�Bc����~���- ..��x�|o�$�B)�b#�@g_+���ғXJxm���y%������(�����v�����@����.)�#4V?rF=�-�?Y��p$N�qBvGi���J���1٭&FW�Y�p�Y�dw�Ii�+ǰ�nJ���~���|6���'����	��o�J1ρ���z.�ZKoy,1v�)L�{S;Yz�
2��T|Զ�9���`�ӪӁ�Ⱦ��9T�UK���T�A��M�8����[�WO�����+�y'�&�Ĵզ�bo漺�` �+5F�8�W��	T�*/L�ŜJ���,��j'=悏��k�P�tՂ�<d��[8]?͞���U�C�0p��0��/0�M�=�6�ِ���M���~a�1���Z�:��w����U:��iLi4�����2%h�CWHt�,i-��%ӻ�N���.%�0ؚ_'�:�9�B78��O�U|Ѭ�ʗ9,,�����g�x�V�8W���u)6��c� ���mZ8o.7H��¹�4E�.(�n� ������Nm`������)�7�-9��$�������f�Mf�6�_���_Wk}�;�O0�Bf��[(��L푢�<���9%,d����ȗ�����X��W��.�����MU���.�7��2΂*����Q)A��]Y��6M>����򁽷��s�"�:�c\���/�e�K"�RUE����O𬙝����[�)h��ϻ.���ޭ?��X��u�=���Ŝ�K�Я��j����,������пV�q(��SjϤ�_��{���K��}RE ���BG�����D��[�j�_�y�w�]%��s���i&]��CT]"3�T\r4��IX�Y1�8?�wD��q�g�,���ż=7AGW_�r�F*�۳�B�7G���?ԃn�ρԄ<⃗q�L���A����i}��Ex?�=I��_(�^3�ws�)ic�mF�Sf��pO(?R�ᶕ��! �XB�h�!�~&�T�d����!C2����9�h��t��r�f�pX�1�N��qӦ[!~���$��>u5}=�v�\l�]���g����	�y)�>mֲ�0