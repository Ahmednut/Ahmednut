XlxV64EB    5762    1400�b'!?(ѩ:��O �TrR����X]���&j���9ҹ������b�d�8��=�[%Ѵ2i� /����,']���N	�h�Ϥ�/��xO@���H��W!<���Q)���:B6 �����{R�q4lv#n�Q�u���?�¥%o�݆%N��_���b�W�	�r�Z�Q�����=�R}��j,i?F�%�֛h�ຕ�&`�8p�)����z�dp22����!Ü���� ��bN�r��&�,̠��9SƟg����E��׽����B�N�������  �=t7����:v������>�)�	@�H˞1F�e��]�& �Ao�����]*�z���wU���;�� ׉~s�o�/yur���&��&2TEļ��8��ȿ{h�X��Z���dg�U�רO���fhA��<��4Q=����ڬ���*�*�)vh�=$��lB밣v�G��Љ�e.�
`�F'��[I�ۗK铵îy�l��X�a��UL[(C7���鴥[8�F|��TnF�IW*��R�ӹ
��*���y�k��AMg)���ٽ����G��l �+b��/XX��D~�h�D$�͖�9��RӋ�~��`~��HxE�����3^�:|�5Tv�t�����OaƊʡ2��[d�	��� ��r>k�����ڠ/�(U.��؝LLa	��'�M\b�c���0�C��TR�Plk�Q�� ���J��d�B0�Lu�!6�t���g:���,o�1װlj��v��Px^�by��Ӥ���j*�^���j9�q��qV`)R->|$r��T����R�ۥ H X-,�1`6����#|�,�hA��~��96�4�pWם�{W�� �̳�E��ӂQ��Ǔ���!f����m�L0?Fj����eS�k��FH�����5�C��,�B����si;�q	gk�i�`�٢}� �:Wm�=�s��Ť?q�S��9�V���'Қ�R�]�VkN�%�:V>���g������`���������\�z`�Ea=rT)��� ��Q�kW&P]��X5:ǫm�S����&u����[YM3+����z��us�De�:1'���)��T���x<�򑻞���R���6ź�|��!������Y$��Ɛ[��
��}����]� aFzsE�'�1	���7�YK��ߴ�mh���FX�8Ҷus��sp�y��n�0���I�9
�#�#�$��e���4�oeYP�!��CU��>�;��Gc���j��Ճ
e��]rolD�"�&0oϯ3H��!:�VD���,4P)b��������[Uk����ׁ!���>M$��'S���ʀ�*u���եЪ=j�8�iC8��|�f��f�]�X	��W���+�����
t���@���6�NpJѧiDy� �ܱ�&��{��t�v��>ຝ�]�$���+j��I�h)�hM���9�ӄ���d�Cb�_��D6p�r�LR+5�l�B³��$��96�&Bk6����D���2FAD	c7��HN�n���{c-����?�O[)�+���M�Gre#v�``n��/���. ㅮX����`A��p^�T�	�e�T-�z���l�i�2Z]��Uo�D����aa���5D ���7Y���YWL�Y�Gz��X�����93��B"~�B��XD�51�K��g�h�������(��A鑴*��3���Ro5cKײ,LA'ޚ6�$23�:<��$��EIJ'HT/Bep��O������fU4o�{(� b��zO��I���(�]`�-]P��#k���
,�Ǵ0�)�g�b�Z��ɡ��Ř�ޭOM�%h��Ng��s�<�X��%�oFfG�psܰ,Qc8�@t��jȠ~��C�/"d��w��D�M�2�5��F�	�A�S����8���/����5�8���2�,A�0�����g��k/%��P�4{����c��R�Z���@k���}̽'�*�ԙ��)��yJ���L��m�E�q&�9��ish��ǎ���	�s��@L��K��B���e�6���*y���@�+����#�`A�=g�RZ"m�����Kz�ĳ�$����YqxH� <I�>K唍tPOf{QK?d��zNX�-i$Мf�@n3J������<�x�K{��9Ւi4�C�Zv�|8����k�9��� /��j����|n״Ae�8�^�� ȷ�
�D)��;��ł�vhw&��Xf �|�X�>x��A�!�2W��~�o9ѯ��흷2[^т���&�{D�㌗����P���z�1�Ho��@Re&��֚���c�y�+O�������rz��.gC$��,�1���"�'�5�0˩�#�)�>?`��#3:;'8<�3g�������b[1��t��Z��]����G�1W�9�����k������6�Ñ�9����+��F
q�'ؖ�a��tI���:�"��8��N��~����:�c�Ͳd>�\xT� )4յ��@�����ܬ�BB'��X#��՗���g���s҆��~-К�q .�9k��^Z�Ί�����o��Ox�A��}$]�[K<1��6�\}�{\^�wrj�Ż-�z��Z�0�R�n{J=��$<hA^ M�����@���P��>z���_���绁��R�wؑ�єA��uu�a
®k���8�x�#�ա\<��h�����k�����|!����l�a.�'��u�'�4��U�Ƴ�:f=GZ�P|�5��_%0E;Ԝ�K�P�Y�]/���8�AR��g ��@�ˈ���	w�TtV�,O�swn���ZX7n���Ϩ��`��a�w&t��	N�W�w|��5\�ݨNG��q���/�L��7�ixPy����@D�<�mfـ�d!j�Gi_$E��&���S�����}#5�w���f��hؑ���{x}�Ѭ&�[N�/���;����B���+�+~��e��	SF����2�s�@�ǘ��^QbfZɁ�Hl!�8]�M�F��E(Z�mkDH�|��:�޷ڒN�ՙ�(�P���6<�䝂���`u���F��,��R�8�5;�%�:V
2��O����8�H�2�|��ѽ����ꮥ�gA]=b"^�����r}j�t��o���G��$�)�('Y��O�{��H�3�����ՇC�/�3Qb�E6��a�,������J�LZ�SN&��Q��Cl�MB(���׮i7���>��o�y��uX"��'��o:��f	�����Z���맚���ޤ����L�&Y�,P���K{J9�m7s�snZ�3��\�����<����0C}��qR��VOUW;��_�3/aD��_���p�?��l�S�_�ӎ�q���ŷ�#�#���j�H�����g*����Q˃E��AɕXz���<�)�Ŗ����F/��K��,2��:��\u:� I��^6Sb��5&!+tu�v�R���D�#ǭ�
�C��-8�g���sw~��?����ess�.����/�"�g;/o�w�S1#��,�T�����6��`������v�{�S�򿓗�^x&m9Y�Ϡ)\*��PI����N5_,^Fǰ�ٸ3]0S��<�CX᏿���� t� �J�e����R;@ILl�Cf��P���-^ڷ��h��~�ɨ�>�;*�T�U�hvy)[�&��� y�mVC�����aשW���M.�cyzI+�"\�Ç�s�@��ON�n��L���Ƞ�.��kp����߃�a���ƒ�7Ĕ2�3B�˿L3���Ͼ�W�
ڪ���,5��-����%���o��}*�r���*��X�.���?YIXذ�Is�Oe��}hY���*z�#zJ�L�q�����8v:��P�):�%��K#��@8��*;�kq<��t��wߐwFʏLɬ
�0�s���!��?h[k#��$�����* ;钻98՝0�;@gօ<;Kov��!�t�wSpB�o���@�t�	]�Z]8��ʨI�2� �e�s=G�����:�׍��`�;g�m[2�d7���W⫆�/��.��mb�I��U�:c�?7�����$i����wP��q�Ok�c"]�{��g�)�3u��hx:F,w8�/w%y��#6�{��jP�,�=@"�FbPÝ���K:��:WU�y�88fˉ�yN��$R�"�
�'�R`�
�[�Ձ�#�����s�PȰ~Ԭ��h�b��+�'��mA|݀��_Xj�ovm�����WD�פ�ؽ�՞ʯ����������Ӈ��}w�Mu}������)*+��_�s� 5�������-����(�7߆��������=?��䛆��7D\[�1�{�� HR���t��6%Ϩ�(�-�o0�1	�(.�B�1�CD����Xj�<Q��#�k������.X���2�~;+Q�������1oN��P����qR+����	���&߻���]���$�;�� ���KL�&F	�7��6;N{S|ـG�Q�P�F�¢��R=���e3�C��jq�
�2��3%�(�)��|,�Z{�,�p���(����b9@ce�m�:紑-���0ά���M�
�j��8Į͙k����y�D2�ܥa� ��s���P��[���!��m�S*������F���ϣ�Ke�yq��.��o-I�ڄ���� ߞ�o�#��s5Ek;�u	�G֦��-��	�ƫf�H��BĠ�&��˨� �'s�d^+��3�Wg-�!⦌C���Az�Z�~�>6.���w�}�¢Xk��)�N�Y?�HM!��p"�ٰ@�ذ����o�����ɣ[�	IXշJ��v��ba�n���n��f]�$>/v!Td��=g�v��^�Q���P���	�Lo�y�gZW��^������b���K��Y{�qvO�$N�#������d�
0����D��B(�ޮ'�4k�P�n�	Ӻ��n���bɂ�*���N+V9.K@5)�-