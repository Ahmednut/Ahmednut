XlxV64EB    5739    14b0I�,ěn�Wbc� �M5�/h��L���������,���Y�';e��GN��47�ŕ3<^��3�[�e����>��V���P���NKۨ�-�K�m(�*���Y6����YX۝��-ho�US��ҋ��
u���:����Q3�G.�����5S��o�EAsyrA��7��5���mz��C(��b��f<׽�~ӯ���
�U�2ی���^*��������ֺ���|�1��TIOr��v_\p�������]C���`|������V�O8�ay\�5JL��g�a��{��
�DJo�m�A��T�C����<l�ܞy�,!A��f�}�y��^T�e����9lͨI�z �E`ǹ�jLh�}hx�,�2�}�u4?���|S�@i��R�U!�.׺��pϏ��j:?�/J��m�I�{�lp"DX��y$Kԕ�}�Ep~� ����-�{4�R������J�9f�O�l�pn?1�������Ơ U�T�8才Л:��;U��9w,�k/1�0�<|�s�dz�O��p"U���|�WA� ��2.9���-�����&7��Ɇ�� ��hԱ���|<�Z���j��wrO�tq�S����3?��}L�"�zx��5F��觤ɹ:]Q%͙q�5��!�$���h�:���j�p��D{�uE��G�w���+�4��V����ڜ}���Vݜ��Ώ{� 
XJp�z�
������P#���@���v�3!'�ـ5X��`��s�n1�Z��W9��ORk�*���[T���\r��yb]K�oDq��v��j��o!Fy�c��i��[��wn�U;Ɠ3�?�,�ImD���.�+����-壌 C�� p�P}>��Nb����82���\�te#��;�UKr6eh}R�V��Y�m6�3���P��"@�&�G��~������^Z}��Fq��S�Ճ�\��=��k�=��짴�2�ME�bd�^fw���NN�=��mHx�A>�P�}w�&���^�PQ,վ�F��#����[S�	�
�Ё�K?۽�*JB��|04�pПG�"�4hK�#����%:�;�O���x5jt���d�."{bʗ#����.���o�(���/����NC�U�7-��\0zu���b7�#�(p��$��W�OW�X`Ka�k����\�F����ײ�3���ɡB�2f�у�=l�Cm��N7���
)�*um��m�濟��ŀ�ϣO��/�d7a3�A?uX��$t1Eb�Z��i�xM����T^��ԑ�:/�/��%�e����2I �*L��S�*�H1�v�=HϖqX%,K ����@Qx�HP%�D/2�w{A|O�̻g��<������	��z����Zw�Ai'�l�'���$�M�O8��WX\`p���=�2��7�נt�� ��$�1|V��������t�
!��$�xºC�IqĀѦ��ޯO9Ǥ�Y��k��;cY����/''wg`�x�����l� �P�Nq�nE�����D���Sh�IU�Tq���a��T�G��9 �b��T�BY?��̈́
��΋m�Ɗi�qL�l4�/-4hI:��~�|_���+��uC����e���O��l��{*�	+���Q}j��jш��y��tQ�r�����q�Ӻ��X��N9!0{.����[�;��ϴz�
�J�����W�N�	��f���h�C֣�P�v�)vuӝ���m�%�E����m)S��hP�9��jbn?��=3B+{��zn�E���] ��Sb��Ä(�u4PA}����
Z�	4o��gU"-p����+4�6�K�Զ�&(�rb<q�3�|��* ��)�
���G�Ծ�oi�6.|4�������c�R#�[�J���ox�G3w�/Y�D�n��'�)��_;<H������@Qh�D�'�9rC�F]�0�C���g{� �n�C+��m��Ae&�W�]��kȚF��Q��Jn��QC�@�ge����Sm��n.�[��	V�*r9�w�{(#W�,��"�ˮ9�I9�m´$&+��a�K;p��P;�������-�P���Ȟ_��C��.e���������ZX����#���$�/mY�~v�z�An˵�]���9 FyN�.	�6�� V������R��]�>��o ?�H�4DT��b�T?��~�]�5���@0N����LNd��3�L�.�\�9 �r �����t�{(g0��|�����}AN���iK�|���&��1"�cqfd�bm�����c��=@	�أ��w3�U��i�l�c�1^� R��2�� �����4AZ���۩W�ӕ_"J��\�F���t�/������<j�_Z݅�. ���A�}�Y"qe��ݣ�#`��9[,�B\���ju��#[S���9��7�1��7Z
�����[�X�ן�)�tCP{�m���Dq ��}[ʑ	�`0+��'YfU�F�<� �S��WqJ�Z[.����ILWtځ���L�QEd�H�s�A��跾�ر�_9��3@8CC��;�I���YH����j ���Ak�������c�J�?룡���K���xr�u���T�:ϟ�=8�+Te�A;�ʺ���O�S&+�mش����H]��?j��ע'@�u!��nU3�`6^��%	=�ӊc�R^Qoz�)[�s��r�6�fK���� ��'ٕp��P[�B��4Ś��J?|$R�t����f<�B�n{ϱ/�O*�azm=z.�h&����>�sA%'�r ���p�ū��`V��4�<�T�@f{����xz�`�Y����J�p�BoS��������|�6S"�����읛�9�����X��6�n�Kj�7D��X
Ί�1���Rm�F��I��w9g�X2�ok84�L�68�kU�������sU�����|��S���DQ=����Eak
����o:�
h�[N���*�b�Y*�I�UO|=�,�b� �@z�w���A^�}�08�ğ����$��<V����E�ۿ�������Z�4��5S�Sm/�'0���ב�0��s�/������V�7�\���(��� lKp���!�4���gR�JI�!�P��x�V�5��wO;�kG�]�����7#��w����i�U|*���z�"��<6�Q�dɦ��;��P��x��]f0�p�vj�hPXc�7��g�E��$j�V�ouG��=b���D7Q�	z,FC��M�K6��t���x�d�D��M�M����ꀅ��fQۻ~�t�-<;#O$~޾��^�����B-:.J+�N��f<sjY(]C@Y�e���Z��E9'e�D�M�Ba*�~�J�2��t�}���h>x���*R���Ô�HT�� 	�8-�b�>tL�/�nI��د����e��
-
��jƫ�J:"Y�U��.�w��/o�?��Zn<T�/L��Px��B�#�������D�� t��	C�͙��m��� �A�y�4ϡ�G#�'�zB9��cv�ſ���'`ÉѶ�M�J��Ӷ�W�P��@>��Ya�n�ӊ�ݧ}g��){�Yk������P̥�q{Q�߁D����������2�����b�
1�^��E���(�~#ܵ��\�`�m�^�w\l<��\7���yu"��m:�cm��:d��0�eο�.�䓀:�J�55�x�c���d���G��X�/f��x�ܬ����KF+�6�{�v������>a�્c�w.�9��h֩~=B����<���,�VͿ2أ�1#�x̶ߢb����%3��z�<B�Y~� ����+x�`U���#�$KJw�E�k6�"�t{ՌTW��N�$�6@�U�LA��!�E��sgD��Ƶ�,p�Q\��X�i�R�$\�S�7�蚖����������E�"����������N��]���{=����#>�m�pr��*�������~r�/��n��p��A����	NE��x��/F��Z��a�gk�ś ��e�.�R�����E+sŮԦf���5�8��p���ݶ2��D���vݳ\��MaX��[�TV��ɾ�CR���QB�[����5�'� �ꡪ���Dp�8@^�0�䣖N#�`�	߂\l[��̷c�%v���.�L��Ը��v�)���P���F���j������~����+��f��/�U%�$r�Ab�w#�9�v뙂2U�2eײ���#%��i�����q	 ��K^�#����t�a^�cRGvg�hHT^�>-`,�3^M�d��s ,=��i�!�Cn�]�h�44dM�݇P�7��#u^mV�'�l*�E;�$.�bo&
�$��R�0 ��6 }#��b���<w�1V�)�� �������4��h�p�$e+�����H�?�(T5�����E�K�A�Aa^��	ϱTl��ZN���Z�=(����e�����6���h}Y>�i��"�dS��>���������'�h�!;���3��9���8`s�%�d�n��I���C���%�DJG����F��s�饤Nਭ�Ҹ�����qA�*z�t>_��gï&���:���a����k�� IioȨ������ky�3�f�����2n{(�y����ħ�?���y8�'�����&D�\�+%���F\����X�W�l��w���&�E���6�ՏÔ��	p�2�\��,��&�/��a��̙�A?j��@	����9cQ��3�6�@?���"�#��ǃ��m����t_;�H��%ͨs�� ��8�RP�e��Q��O����.��]�'Y�
�%.��lO�V�+%P�x肀����67F0���6�lXMR�(�� �P���I-��Ǖ)�9}c���ɺf-B�|7'�W5Q\��o=y�#pO��AV�<mK�=�M"����&�x�M���3�ˋ#�_M�2�6��^�����l��цP�"�4��� ��{���过h�|֊�ҾP`�sЃ�>�w���]��)�[a��C$�r�ք�¥�����巔��lj-#k�ƺ�$(�oN��j�~6�{#�Q�w���9��L����k|��'M�	xxE�/�V8��?A�3q���ሧ�9����:���)�K�5k��C҆�
=��ْ=��֚��(V>������HXLE��R