XlxV64EB    a7af    1bd0�v>Y��.j`?�ͩ��K!�2�������,�+ǣ��"�1�l&�RP_�$>s#f���y{��a�ӫ�zە_�]&]�m;�4�������ug�Qg��ZR��$mI %�(�	, �mY�O`7�R4�LA��.�\�7�r���؜��3Z���3�'�����UbN�g�+~B�T"�Њ��a��>D��H����!eCmH��GQ��:���+y��o�J���`�̭'�/��N7�vx��zrP�l�P%��}E~�r���en�^`+Ǌ��c�M�W�G³�3C\�I�٣���Z��kb�%O� ayh�?)�R��J���P"�2��f�ׄB����B�K�+S��j�i����?�WS�������Z
�8��m4
�+�5gIh�*�&�#k#�{(�P6���8vc.���k�{n7��� ��9�ΗX�0�wmƠ��W�R�l�uz�"���`I�dW�`�pzr_�� ��J�UN�g:bhE.H"�����>#�/3'�bw�kB	i����L�2���ݽg�������ׅB���,��iSs�h7�y�%p������?���y�L��~f|�g�zҨ�Ƈېs���Z%�*����c�����1�@v~[a�XbyEe���|�?hM�~]��%�~����" ��➳�Z�Gl�#`i�v��J��l���0j)9�~z�o�
Ԥ=�s�_Ĳ��sߚ0��I
����W��<�i�#B����N��R{��3�ny%K�%xB�!�_��@ӣ#���p���2���}"LN��Mt���]dm(��(5�H�<�ݸ������nx�Ñq�OL��C}Oٙ���>�<q��Q�x|oL���G?����|��H�������ꁭ���֢�jjG��U]�)Egw���j>�ʖ�P5�p]A.�L�/�l]n�ɚp�t���� ���=��t%F�Vۖ^g�
pȁ��
Z��7'��� n��~�I��=�=K���zu��CM	$34�ߦT8=
��>�<d@���˖ɺ�] ;�t��IB�����+��R]�Z����ʡ+k�Wc誳�٦Q��n�@��g�W�3��H2dVQO� g�8�6��� ֣^�ȥS[�-De�x�*�Ҷ��쿅�k��������f6��_��GY��;��0x/����Zd:�����u�e ��.��IR�w ��pǧ�lׂ̃T�NB��jc����
m��&.�X�#v.=�1,u���w���.�󏪱���tN������aW�h���N�)=�t�Ш0���Q�����O��\�1wo+J*>��!��d���YDC\R��$�E��|�vJ)w����47H@����������Om�̽���X���%�}h�nbحRw�ǆ$>m���2G���E�:��"�.y��	e�8���P��wo$�7 �Ձw�lkzO����� ��٭񟎨��b=��B�hy5��$����š�O�O��պ*6.ovf����d��al����@�)�L���f�,��˺�N��OOˮW;��@�%��j��n�>o�p�Ċ�Դ1��aiF	:b�Kd�	�(ޭe5OWJ\`�d�{��M�Y�N���Q'2�ı�Q��0I_��U6�Nq�b�4}�W���}�޺`���!�5�(�M�?���J�Y�B�CN�,M��S�728��v7�?��6�v���5����aͤ��ö�_b/�xê ��X�b�ElޭR��vOr
�b�Ic���wC�Ł�[-�pɅ�dQ�վ���t��V�TF�LDe_Cx؍fI�L��w�t.[��b�i�x����8!�2��C�	��s��P��捹ٕ"2�:��(�{|۬���k���k��<t+2cyu�C]}���Z$�M��5$����.�Q(��~ʆ�(N2�r��3�����3�O�4�D@����V�d/D�f<��i5��a01������x�ԫ̛:�&������V�c�б�'�;�F��i�����&M6��e�B��eIW�����4��MS�C���؟�:�tO`o�ګ]�N	����0��4�D�|(ǂl�Q������*ϯUcɱf ��}���V����s��]|��$�_�4D�8��I���w�-܅&�JE(��z����q����i������XϮ 9�Q�yޜ�3�����^_n��
*ߒ���;dg�)-�/�
4��U�:�?���̱��"�w�6gע��h�O�v{����%MY3;\o�L�* ��ƛ����:��FS�����"x:�����x(�cg�l=�U�sG�����DمQ��@�� }��}��]SF�����	-���S/��4�����rƚ�8���yy24]�u��P��7aд����3��P�4u�i_!e\���H������l��_�<29f�)�`�`��:��o6�����u��ͮ䓍�t�G�*�N��m�NYC�$��O$X�4�!�|��@��)Xo���gt�������I�ll�U�$� ��go�Hp���jt~�څ���a��+�л+> 0fj�;]��3;#�lI��51l@e�?ts%g|�SR�Z�j��ɢ/!�Dm_*�éY�>�rG�1#_��:t��r'�V��Bܢe	���t��R��L�*�~�r[jh�K��_D! ���h\��?����>�u�.�&�p� �p]��Ao����1�B9��;�t�R�2��B��&u�h8p!���Fڍ˩P�E�Ôb!ސ����z!�}��f[Fm�9C#-���T�l���0�*���<ٮ�8�L�V[y�W;�K\�o�Z���ؐ2!�]j-�''u�f���bN6X�Y"�����~9Uٳ2l�e�S��䔵�>w���l\�ߘ��sQ�]�ǣ1�A'B#�k�w(�M�]�f�Jjmθ�	S-g%sM��NZ��X����GJ���Y�!�i�=h�ә>�d?�����2*[���:��2{sg�P*�yt~������}����i�$��R�|������T�q�*	r2�/<����pr�4m�ds�c�L0���_�]�8��^D;FٳNO�6��]��!^�^��rY��Q
������H*�P[�j����:��H\øz��aC�nw
'7:�띕@X��C ����r��	�ᓍnM}Oj4ZI*$xɑ�J�E�hd>g� &�mcgr(2��j8L�#�k ��8��S���ޥ~�@�qGYI9��	T�{��T��w}�͟'�=���P���֙�{�/'rv�1�pC!�_LQ�k@�j�}���R�A����4B0���8}?b |9�0�-����XTа�R�Dܻ�k�ģ\�����T�'���Բq��/�<Z�|	�^�z��3n
E���C�������|1���� �
6�^�J�0F*eV>��6l��R������l��[%����d��ΎpA���!�^垘�>S��b���؏���cPHY�}Cײ@;��?"_v�i�7�i\:�������Ϋf��8���@�\ Z�tv�&�#���Q��ܞ�F�-�%T�%�<}��s@G8n:�)����e� ��[
����"PUm����P����B2IוW=�K}�8�Ћh�4>z�#C���*���Q���<T(b��-l�[�&(@>j���Ui
�^�c3��<5�A���n_��w�з�!���˸p�$s�~�\%�����P3�����z���7����U��� ׇ��ӦK�@Ö�����6
�=Bq�S�C[��w����?Q4���٭�R,'�\�����\���u����O��v�F�"��xG/K��yԺ:�R%J�Y�HאI��eұ}�1�f���8�T��;l�ON�FЄ��{�y�Z�-���D\E�`�]o��ۃ��X؈I/�o���e��N�x��6���Q��wD�h�u�͎v+w�L�M���}����n�<%\�
�V��پ�tJL��Ӫ����?~�l��^�8V,�ɀ� ��}�Pv�}� �=j�k�C8��a�8̓eR�Կ��X���c/h�w&)�U%M�|��*��e�ճ���Պ��P����s��7�q3� ��>?�Ze2�Yw�ꭀϲ�e`��!rȹ��9G���P$ ������+���^� #�t��8̃s��s|�^�Z�c��9�k%�����6ZH��j��@)8Y�15�,qr��e�E���� j9�Z2�*)T鵉�!�@�u�.)��������mu5�]��b����Ƌ�L4��V��(�}�t�Ҩ[W#
TM��-�!�5n���J�J>�TK;" NKk�R�x�1ܿ��!��M�$��_���ɈT�~�Lun��h*�'&�]�#+��� ���Y��N5�V���)z�ޯv<�$�̈́n��>����^�1��)�*+UK�ڈV�]���L������9���p�7|P�4�g�2��kS��TU9��Ňk� vwR�|i������1���$)�����^�2%��U��P3<�PČ10x;T��8�P�Ú�<X�=w"%���ʡ��Jn Z �n��+x�>�
 �!�1����=���EOj���̅��0�u�N���J���fq"��ޅE �u�����D��O�0j˄7���|�<���6<�$x]���5Ի���JW����6])͒��Ȁ4}/7J��7�u��I����;�l鋇#�n�,�Z�|uo�n�I�� S�z�|���!X�y�EV~��G�'�ԅ�Ds**��j���A�.AO��E�D��W�d��1��ٝOi���)����{w����"H�_i����":o�Q�ZΛT�����G1襁���x�����`��zb���AO�O�l~���䦄�DZ�)U�ǋ�������F��/ٱKj<�WK�%)[Ǚ��s�����-�T����L����b(O94��s�,�^�s�q��O��U�_��I3dz6l���B����p�x��0��;&X�pÝs���L��tT�b�t��L2�
l���Ω
X�,�� A�����M�F�j9���"�P��*$H�K12ud�lX 	�c���1ULu�S7m�FrWl��j$+I�����Gߙ��}?�d1wǹJh�\������W
t��I@R��Yg�*պOH\0)��Ap#��橳S��CG����+|@��<,j�݊"�X#�`��<8{}���`a��s�;��\��@;���i��5u�za��V��qP��Z$&�.;��ʉ��蒬��گ�׾?�p�/E��X3����(ֈ[Ma��~��Oܵ@e�Kg�PԲ������}�I�t���Y��Eu����� ��K7$��[s t��8N���_��o(գM7j�$�eę�Le���_� (=[x��6�Ó�n�p����ۆ ?>�8��Y��8�$��̦P�w�;6.�̡]`,z�ޠ[+�YW�� ��:�Z@�����r�^�����_�	'GAXT��-��ު:%n�:>�K(C�zd)�m&��dj$�|ٶ��R�-nA�R)t�������w߼'i��h�2���p XB���7��.���]$�ӡW�ퟱ���"�o�A��0��h])'q��E�C�8^S� �vr=��熴�`r�~�Q���̙�>c�M<�Rb|/9y�����X�Z�~�K�v�����z��hҨT2���y;zF�܇��89���(u�@�f��@�6M��Rn.���]Y�z�9G5ms�S͚ "���)y@.��~�5LσMt2����9���ߦ��l#@D����$���v	0�ub�c;-��f��%��0�,q������W��(��z�ͧ��آ��Tk��N�Y�܅Kik��~*ݷ�9#^㩮�ʅ$��=�$ڹT	�i+}n�cA�j��S�鯢(���B�ݼpJކ����o8��Y�����Aj|{+|̨l��M��|i/���;bY`��6�<J�'����`83j֭-;Lo�Z0��O�R_�p�l���q)�v�<���O�ҭ�yz4�/��LZŤ|Ǥr�W09�*�R�D+R�d�.�Ѻڇ�ť��תtH[��~e�#��i�~C&��q�txF�f�*���Ja>WH�d��u^�+�^(=�x 	�4���ac0����!����>�����wi�
�Zh{G�R���@�z�\K<Y�r���`&#���y���M9r��G����4��]O}��2�BNK��0f��%��	��\B�z%~�3�:W�5��y_^��E"���=Y3�2H��9���J�I<:��.��4�����W���W
�����|���Օ:���Hk��#����:y:O��x!8_�,*C2h,� '0�zgp��"$��k�i�;!	��$��*�cQ+gP˺�����>6������,F(垴
m�f*�3�E���ސ����T��a�����j�|��S�TV��o�`�=�i1��O�r��Y�]=��XC��nL�j�m��;KD��rj�����)<N�so���K`fyu��\�cm����f��wPF?�0�p-kr�Q�Ef�TL�u����?Pq~�qS�F-�C|<D�mW!�ڷ<�	+��G�N���d��D#&ҙ3�fl)���O����Vg�/����R{����y��2l��Q}��#H��3\�[�)�����`[�?q0���bӀm���i�� �~.����Ն������gŲ��̶��Ӣ�����.����i�َ�ҍ���n�P#��-�H��\�+F7�:���s�=�~���۔�.bC��E+���ؚ0��b$lַ/c-�`F������o�:����^�Dhc�?�ֻ͸MEz���:g|�aV�5��A�gEUr�6����T
�r
����$����\=�wL�!��ӓp�����|�Ic#�t���o��e�+$���hI��A`2]PV7��ELR^\&���/�Pi��DU���2�S�'ʭ/?��䖖�����;�Mx^4��#8�r�)t���O