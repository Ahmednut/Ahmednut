XlxV64EB    17f2     9b0��b�O�� ��z��(�L��]�I��������+!Ƿӊ���JTL�� B��4�u٣��5dW'o(���7���v&�LU�`�yY��LL=M��|��YN<(
�n�<:W��R���Q��y��^L�i�2�o��q��?�2����q��bq��C��#��f��Q�<Wg����T/,��	��0Ð�h��9��z�U?I�������B-C��%^��������r�I���á��`Wh�_�\x�m�����1�G����Vn쮧%�w>/b�dж�D�ڶB-4.����ψ	���g���Y���^E����w,c=sG�=�X�Bp"����X�s@4(�;؎�ZI5���K���VȆ�^ѥ����Yw�-���n�U�i�jFL*`r̵Ǽ����������_��\1_Â[�/.��9~ўC�٥��*�$�ex�[��w���Uq		�
�?�ou����L�;�E�!,k�!C� �*HD�㻫�}h'q0�z�M[�#�����hi�Tx��.�;���*/���� Ip�5C
�Əә���~�x��Y�Gz5E��e@8L�!��l�\	�y�k�;�
��]p��~$�~��Q]�B�D[W)��eV��X��&�20�ɪfD���&g��oݭwy��	�i#|�>�0��wx�9n��N�zs"F���*�ɳG���Ө>�*M���
9�2�D.^-�	`���TxtQ[�������ß���"��>�:y�)ml��}�܏�6�O�����,��p}�,�u�2���|��1� <.eu#E���l&�A��w,�H�E��6���`�:��U���i�t�Sء�"p�T�BqS��wP�����j"C��N���$~d�ϑ��jlC��yH��1LL`@���(�ǞƬ���+��� �]#W�'w}�f�����$�G� )�#m�����X�+>7e"D1���q.6C��d�SKJA�Ͳa��y���Q�/�U�P�0�;S�epL�c>�.�W�U����X�`���'��|���vf���rc!E;�>�GB����]ǔ�u�@ �����A%�;��M�""�<���B"֘(C���`,/X�=��t+uZ �dd�I?�e�ޞ.��qir��J���3���r�t�k7[��ʛ|�C&��l�� t^,�������v���\�������b�'�]l$j݈�O�fc�_E�t���l%������Z�
����$�����ghw�tu��:Q��}���G�\�D���q��@��.(��Rlb%�V���.{�d����C;"A�S�z� @�Sl��̔�c�W$��ؿ��j��Oj��h��E��@�����G5ä��a>RM�3�8 �F�˟wQ^���wmT�)V�ua�r�x�[d�J���/$�(<� #7sԲ�7�Q�ƈk�R:p����l?+�\�H�憓�$����-�a=Jw��c��!��;� ,\ �M9�E�� ���_�KM�+�u��T��3�o�����b�%��|�
!�����dB�1=ES��e1�%�΄��#
��C,J�*�Zr�0�]���-oR���7�]��6�׳'o>��v�z��u1��8;�[�Mי��{^�o�tI�Y��5)hr�;k��8O�ɟ�
�L�H\��6�t�
�Q*�0~��w5�J	A�@��������/8��sA0�M���1H'G��y[�`�H:I�=0���������F��7��jo*�<9�o��d�Y��(H�9]���?
�W�v�U�[*P̈1�M�qIA0�[�'��n�AT���+.]ե��5i���O��������E?�͋lz	N	���q��i]�' ��S��S�����ruu6&1md�Ҿdת<��Qw�m���CL���c5��$%.���-��PK��]Հ=3����)Z8r��c�l�:AlV��z��ʱ��C�M�E��	�x1bB�؟��%@�Sw���4����k ����=�]���1\�1�� �������SdF�_��֥�����^I?ļ)���Րg�ӓ�`�-.i�7���V0��m��ųvmOb�Y+?���	�ѱ_��U��i�2q�r�`��Y�=r=�_�^�"�����=�` �f��	��g��1W��E�]�j�m��E�����-Y2�M�8!y%��[g�x�7�W:f���p&O���͉���_�켱wx/5�$W:�V���8}D�@��݌2(8�v�8qt��H�	���ٲ��hD�r��q�}�ދL�e�C����T�]2��N:+�#�=9��ό���odG+ Gݼ�jt��X��8EC�=�XbXP�I���2���7�R�kA�q�X�u��&�]GM6�E��A�}q��О�
,T��j���p#L�fT���;\�>�����f�k1��Fk