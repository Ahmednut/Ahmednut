XlxV64EB    243f     be0&���%�Ċ7��qe�T�TM-z-��0������/��?�r)u16��%$g=lD�9׻om�,Z�K�-�Q��`��yԝGhI��A��E��5���U�-�F�T���
tbo�KV��m�r�R��l��p7K���SOlb�9��9��Q�����#ʲg��!�����JS��u.Igҽ���@�+	��A�H�B��K(��-�C����\/I����k&"t۫�,.�HD�	��7��]M��T���&�{d��/�Z$=�W�����t�����5�Dp��Zx&�� |n��WV����y`�Yza��yݘ5E~l�޶V5wB�2�]�Ο�J�l�n��ht�T+�'V4.������4*��!>�.���8i7r>�xۊ������/�m�yj
/� +�������)�_>X�d&�>ox[X@�p��sK��3�k��s���4>�Ng.v/t�=ܿ���2��cP �~��iC�o"6PI4M��ﺨr#�~���ڗ=uY�U$L6Z���i!ٻ	��e��N&���,�����!��y/\��^���eJ���'���(v���:�E��F�h�yOH�J88˻�f�#5�Hu�B..w�"���.�"Ih�9tbD	nY��	�ŀr�v@6�ѷ�o�a#F"($�Y�i8��V�n�oX������5���~>h�Ւ)�X9�l���s��r9�]W���-��G Wm�}�)�1��5�[:&����FZH�%̨��+�jB��+���0�^�I:H)j��
wΜMӔ#>G Hx��Ղp����j\��[#N%N���Ml�t}��N�L)�o���p;�9���Qpl���&�ُ��_����Y	o�T9���#�Et��EK�����s+�<�v��Ș��p^��%��;��I�a	����]O���w�4�& #��v�Ď�Q�3���$I+�[���d�e�"RO��tt�8B���UY��#�����~*���*�~�Xa^xl���,���|�[���<{����4W�O��:�Ss$P~��(S���s�=�[ �M_!36wѶ��0Q��^���s�٫�V$L�	W�,)�z���@�kd���䦭�
t��G"�d�ܣ��kwm�����.2�ȩay����q���F�b�
|�s���ē�n�:���m�Il;WǼ�3GĵG�� j#��ف=`��M,!i��es�F٠�S�_�������aN�^$�b�sJ������3@���h �|i����{c���.����+u%>jxe��@���w7���8�U]���N!�'c�R
Wl��)�	qO�L6h�X�`[�:q����Ձ�]��V�N�?��a`<��a��z�r������nv�h�����0d�6z��"4�!G�F ����5�<sW��oU 
AҒuŧj/�,�6��].x,ɒ,N|�P��s����V.���x�QO�����dR��u�������`3x�܌�d�WLai�%���G��5e>�<�D`Y�k��3�󙚵kF�tf�r)���� [6n�:�a"k77aW�h>�=�a�i�ސmd|�[���r�285ѹ�m���+�LK�����gm��5�uVHP2�T3y�5���ٖ���͟g4[��T*��^e1���G�EX
�U�p����0u�F�u��G@va3��qUĦq!����Ԗ~DF����ҝLs�ȇ����<|���<X+�r��Gp�|���>�2���w:Я���<����%��s_������������C���q�`������b���#A옻�@�ߑ[�����i?�V	Ӹ�Mz{?�̋h��_6�l����G�_��ٲO����T��O��]{�&	�����;�f��j�"9�5����l��5O��X��mGdam�uһ%4f��E��.����!8�|�e�.W��xeT�0�,�%��b�i�j�x�e���+K���">ׂ����eZ���$ J=�R�@�	�.�Ca8��&���b\�L�k!��)-;��GfH&;"Z����8�w'%�9HQ��P5��p��I:UgS��#mX�Lt*�����Ju�.ɍ��S��y�\pvMƻ�ݓ�$\qw��'��#4k`�� DqW��J�4�q��Z��uc��r��	��G�� ���G�һ��J�g�����A��ª��6��N�G3g���Id�܉?��/��M��+b��ɏ�u7t��D�k�g�,8�#�y&{TA��������M�Do�S+-�w����Հ	�+�*��8?MM��}�$�K��܌�F��wJ����T������J�F	�ΰ=��Fԕ��#)&k�U:!�t"�&�E��y-4Зj�D_�����wgt�=�%�Sd��T�c�%t �?�DH��Ƙ���k����EƹU2�0�'�!���c\��^�r�kF1[3���+�ܤIc�&�n\���Iɲ5����0n�:�֖hx�"tZa-�D|j����m��M�w���i��%����vؼ�nõ�����(a*�8��k/�ڌ�6Ƴ���s��V�JE^Ӄ�^s>6�3����:�H���ˊO�:�4~��%�����ء�WY2��9��2h!� {t�撗g\���<�:J�ɤ=[v]�h��d��{l�#&.�����+2��E�&�a���U9W_G��	��~����(� ��L��* �L5K��h�+&i�[�3#�ڎL����N��g�I�ǲ�o��o?��X[W߷��������G���6me�@�*c�a�\NJ���jD+ٻ�q|��8�i@�v�*5�C���,�e��r�fL��J����u�������#���ڐW�+$���_�W��Vi�
�E��	=qyI#��ko$k�ڀ���;�YN�K4=�M��W�>J�W��"�3�3��ܫ*(֏�Ȟr����p�����S9����Dg�3T6ji*�&b-m����=ޠ;�UYd�t�<���N�`