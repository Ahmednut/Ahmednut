XlxV64EB    18cc     8f01(q4ɢ�Z$#�=ʡl���GA�-�e6yg"Y��̣�;� ܭ�e��S���2̪�~C�;��?�.@���8G�������s�Ӄ��y�әc�Z����9��îЫ�Ϗۺ�;zdZ&ߋ�����k}m+k��񟆇-T����9�Y/���g'���dp4z�MF�K�M�Vw��+���,+���K�Qz����]
�rPM��N�&�Ю�b�q� ��{�l۞Rڡ�;�M/K�9�%P�R�N2��8
��i��i���	���xo7,)	}(�yp�'
�-�&��_t����R1ؘ�~k���������ȏY�"�+���Juim�s�ɓA�W�zMqE���w�q�U����=�Y����+�R@��!�;U�PZ����1���):��-�+c�l}f;5N�dI�z=��Ȳ�P�E��W�7��]���+e��9���5�Eo��C��!�V�6O�^}
���/��>�(�����=vwM��م��K����yK&��"j��IX:o���1L:��(��M���q��/��1pkY`	��׏�8����n���r��X9�X�����q��޾U�}���}&��WAgPl�/�kZ��v��
&����`�ν�z<2���3-L,�z���"h��(���I[�y�Ӷ��{��0���Kײ���abQ���:֊�N����0��r����\�/��V�(��/cr�s|�A� ���V&�F�吜ŹPb}��Y��+ю@M�5P�e膧XA��0S�~��/`ޑv[)#������k&۩\񑜿���0��y���ӬNns,�I+�%�
N�+��|0��Ȭ$��|����2P�
�Fz�p4ځ�-�G�k�h6	*�q�����R��H��t[.L��� y�"�Eg8xb%�A�/Ɓ
�F�h��`��@��&1_1a<"<��ֈ��d�&ގ}��$Ӻ9`i��직/� �naM�ݣ�^A��7��H{$Gq��dv�S1l��0ʼo�)���f�jtR~9���]%�@�tG�c�_�}b�N��.�k�s���݈�d��G��
K���-�y�����_�Ns��!�Q�9@�����QZ��^Č�� "�c�^J����զ��G�6e
]i�is|QV6j�������]���=p������kY����̓��S�(�D�A�)8��ӳ/�o�eB{<�$�ib�ceF{��?��]� ��\�tD����ǉ*7H�;��_��lg�0��H��JD�B_ c�HBV9wGw��#V�N/yjn����K=�b����$Z���	�<���M�s�7��VV~u��-`����� ĭ�3�����UnI���?B�L�uF�([��&�xC��W�b��K��v���!�;�vjՈP*w������b*�\-F���'3��3�����:�L�'�ݾ�ƿ�I�.�8�3U��߹�/N�7�1������.��/]��J��������1���{cG��R��U~�a�ZF�M�h�7#��a��>�@rO@�`w�Ȕ�����thp_'G��@l�֝r� �_�;�U���EP��d
�N"N��5����}۴�')�nn��v�ߣH�O?DP�_I�ԧ��y�<�csKw2|"طv��w�d妏A��d�
M2�F�
��|�R�ai;^!pw��Ft�|�-�2/��@� ^��:rq��� �|d�X�S�u�p�~i�B�_��a���N��R=��~.ҫ����q<�k����E�����/�FaO]����?)␙�sP��o-�k`��3�4��D^���ES��u~�Xi�w�oR(.���b��	�A�_����� ����u'w3�l����u�W�pLS������k��1nLUY���5����h%�94��E�X�3I����g����'I��QP�}֨����4D�|h)�Q����SNPeP�^BD�4���Ŧs|��Xf%�SL>��~	�iْ�5���v�9���S+�5�;��
S�<
$Q��Xr���x��q�O�]j*�8md�?.��;{ffN��!�4`X��$�3��%*֡U�Y(8lL�Y�:���֗�Lv��.�׭El��,B`�
�B�>B����O��m3z����|���NJj�7�3Z�����B[*�#\�o������u���G���w�m`�ڦ����0+�ڎ�;��L���u����ָ�H�#{Lg�