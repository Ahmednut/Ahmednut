XlxV64EB    1595     840%��a�@�?dj�d��P�6���w�q������Y�)��������Ɔ���}������<�����bH�6!L�"�W��3�F+���l���@8�s����L"*dg%��Y�U���Fy�Rxv.���� �����2�"�������L��)��,q��Z�y§[H �:	����)g5إx|���>��M��Ik�&������}�$$�yzL׍W�=�Y)�_Bu2�w�m$�[3��t�+��U��L���Z�������_��ʕw�tm���������Z�+1:�*0#�R�J��qi��^g�0�d$=�U6��iю������us�T�_�M;F����DdW ��)���i�Z�)Yh�J�6����1w22o�B�v/\[�C��(�9ңZ��Kt<��e���o��3����g�~�v9�V������<�#I;�*F�k���E�%��z0�@�Wn���>F9�o�* ���� ��/���;�|�J���E���C�9{%`���z�d�>�;.�˹1��ƛ�@�z݅����,�Ɨ�⸊�`�5W�uJ�5k��ڀ'[���� V��{ROo�EA������gLC�6-�~���Ҳ��$�f��mK%��AЄ5���ܰ ��X�CV��&5�|�4FT��5_�No���[�;���s8f}yR�svg�����O�-�F/)��m�D���.8�#�������Оd�6�!�g43y�Ͱ���Iފ�g�96c
�x1%����>r�ܤy��m�V>�j|�x7�K���An�|8�>�tU�oS��1�ӧ��)
)-��84 ��tO(@�U^%^L�NM����s�k��I�c-&�m5O9c�[�3�F8�+m���=�ޖr���dV_��,�du�����E�ET�*�d6�@�sҁ�M���,$����#��j&��g�T!��Ew�er�ݷ���]9I(�s���:��T�8�C�h����Tٙ ����;�nY�~��~P-���4�+����n�=�NEb��Z}ݹ�4�[�eT�hԐ��V���ɝ��޳j�gr��0&�p�J>|�X'=�����#��c��^������'@��E�im��Bכ��w���Oc��Z�o±*5�N����,=E��nϾM�7Z���d�j����������K��qys��/T.4e4��<3dO�ac���
�.l;P$	Fi�H�d���U�B�l���B"\�5ƀȥ�k�m�
�ti�[��j�$qԲ����]p�u0bGb�� X�F�����*��^Ɗ�ZIXD6x�G��LkQ��;(j�$s�m4G��3�Ҏ��&j���f��M�<;�?���1��������P']i
D�y$5`+��AC���V�SrITo�jC�<�d���́�R[�}�IK�����֖ )뛣�J�oi]�p��!.b�Jo*��dS�UAX\�s���	��["��2%�����"4c��`��V��a�r
�m������+�I�Q�'�d�P���-�o`��!���X�x�X����$�,O�V���6�ZF�o�7Y��W�D�BiE��^��F�iOn���7�ם���,�KDPItH	��y��C���<��'�f��!�]~��<U	��+t<��2lK^��$Z^�upFry�qs�Y��1A8��´pZ��v��b���)�6��K�~5c*��	
�,�ѐ���%CĮx1����J��R��aN��5hy���e��8��mX�ʘi��V���k��T�J�f�5]���R��p �0G"�qz\�5�l��#=d��d:�H�L{�T%������5���]�����Tξn���J^����[�A��Z��#ߴ�\e��d.��T2��è�}JUY�{�;�����pq��w������~@<o��B�N�C%ʹ��RO=��%}���YY���s�GmY�����zP�%�kGX<E�� &�pn��x��Ćuֿvx:���'����������nv�ߦl.�["�X0=�Zt7����b6�+�/۫�M'�ґ�a��1�� 7aS�;�7�