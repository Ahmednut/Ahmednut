XlxV64EB    2b55     c40�x�Wݗ�^x���#F
ƀ���ʜ���8�ߠ� �ˀ�%"0�gb̍�z�)�	&Ԛ8}kM���[^�ƺV���!<�^�ƺ��;)h����|���*<zwH0�Y*��곏f:��T��"�WA�0G�7�{U�|��N��7���)c�-�-aO��{�Dy��<N�X;u��4�kspַSd�/Qp�'���s��p��V�=Oz�G��G����5�wʏΠ]��G�vץ�'�[od�N�S�9"�� S��⧾����>�y^��d�qЎ�N��cP�Isw?��g�F�-�G��%��n� �6��s>�p���!��<J,�%9=�MB���ϳ�����d�K�e��,��h�iw��L&��o0�Ύ��G�z����$���Qp�V��n��/AP\Yx�E)׿XQC�L��iB�V�	o�U(�v1;~�i4.2?p ��ե}^��PG��7�̕+m���юd��9�6�d�q���pz��p��bG����d�ڗ"e]�3���m��$�Qᙶjm�����Y���#��Q�U��$��1��#V�7:~
ǈS�RC#>K� �d㯟�n��
m��`�eШ����;[*��g�{�g���h��_ֵ�V��J�pX��aXV����?�A���8<�����X( d�����`�����v.8� f�ʰѷ}M�M�t�sT�e��
�Ԏ�4�>W$�\7���5�r��4ԕ�A�G�Cj�N�vD�&L=okw�!l�y�!`k:^�Z�P7hmmJ]<H��
��\]C��*���K�N�� M����t����~j���	HVs��w�/v��j���/N��a<�B��u3����2\��'�M��{C���T��?��t+���k[Cֻ��0��-�\��V�[Yh�+�ʈ�k��3F���a��������vg����������'���N8&��@��X��*/撯]�S#hm-�����}���0z��XƁ�K�4���L���?�^]��ޟz���L�F8>�r>Ң�\ߜ�����(����k��@&��Z�3-f&�u3�J�	�?<F{���Ңs��|��RB��eC�$"�I��)I	��@�O��'id�B����@��@	�r�X6&���5}hu�<b��t!z9~w���Ҿ��������_��?a	}��h��A4�sO�"j�2ڻ����&��'��A�
�|���)��u�u�p�3f�m%$o(&��S�8��G�q?�]κ[��p^���.Dx��O�mS��X?���e�t���a�c���Kt��V�{�:�6��w`��QԶ��z���iҀ�曊�τ������?�BĜ�|u�T�k�ӗ��:������`U�\��D?]o/XU	�3c0��x�Jt˔&Jx���&;J�[q1#����A�W`%V����4�
�	�#@%��x�ή�s����0�C�v���Ֆ8���>C��o ɒ�_�@�~����UG1��x�ȼ��#�
𣺬�9�;)�MîJtSèS^�S��u�������k_hg����2��w�z3Q$4�� �ŀ�7{��'^Y�P��d����T\���y�Ҋ� c�ș.GfgR��"�*+��>�Ub���2<�7�˄Q�Y}_Ԙ�oA��ǈ_֦��P@�-}\�a��h����u�c���I��u��F�����*w�����r�)��U9�ۗ�p1�[��_�$�BXU�备`7�5��o�ӌ�)'Wݒ&(���W�p��sS2L�e�F�E�m�i���t4E��:�D5ɷ�;�T�.wn���f��~>�10���K	�o��1Z�F$JZoG���6�dو�SC��,�{���]�Nz1���!�g��0�#�bJ��H�j��������"�\3	�5?�i�����mV��著�r�Ngb�'!*�1I($�c��)�\#�ޛ�b���uG�W	���^z��jax��ЬWoY�t���#/����]���}��{C��pb
��R�aT��U�.�ʜA�:&B�}�������ڗ��|�7 ,��&��f�wǖtzBǸ�+�la��i����e���P��sy����I�|�m�tyy/
P�)�W@��di���y)�)e�V|=*鯋3WL{
oN\l���,h���@	�w�3�8N?�12$�a��]�*�_	�4��j�P�q���<�1ԶCh���p���
�F�G3#!��%�L�{� �Z��^��_o:���,�m��"y��s���=^c|q$7�e�|�A�jo�I̹A��e�81YW��S4���8��w�1 D��9��B��XP5� �f)���{������rԉ�G'��t#�+C��g�n�Wl�MZ]x&=n;��IY���Tn4���-n�+t4��&�|5����M��-O��������gl�����Se�h�y��dUْ�澵��K��=��Z�A�Ϩ��[����_��̼�����w��H��!
ۦ�1X�sN&"*e?�KqgLP_\��T	�k��Z�W6��	�K��Z�F֪���T$]��dU�lg�3<@yb�Q���y�]UeMo���S��^�U�y�G�� ?��}lx��Ж���Hb/��b�:����D<����^P=ZS�CϿ�������+�6;��!�.n�� �$�Pb�A�%� ����k��P�gW�V������i[��V���Jj��F�Ğ���F��'�I�G��(��5����k���S����~��B8xY\�[�VT�����q�(�C�0鋽I�N�/-��Ó/��z�w<�[e/Ú�jQ~�h�zS�]�o���f�dU`�kt|�����4*U%ݵ�l�U��|�68 	�O�Uj� ��.�d#�^�C����"��~���Jv���tVf��>f	����k��WPog퓦��3� M�5���[A�o`A�g���b(i� ~�NP��VQTp.-6s����o�;Vz���+�6�i�3�7�<NLv%>��5��ec�XM�,���_c�ɥ�ߙu�.�d`7/�?b����oQ�g��h <���LG�+�%�7���n�`S�V1�a!$����	$t���q�����P��