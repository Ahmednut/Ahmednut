XlxV64EB    27d2     c40�_'k]�О�9F줒�tg��F�X(<�І`y�����!���:�60Wߌ�ː�J9����<�/�
禪�������{����$�� �]�sZ��y`�HG�@����`<��=��=i��D9I���ҹWb�U|T
Ը�1���)|t����P�U�c����C�-��]�YQ��m�ł���ן�5=#.��0��K&R���ޏx��HO1JXϳ-����%�>|xF�>�<�K�p�g�Z�<���"^SWo_�:�� e&�kzˉq#|��}�5*�h���>��87����+��)�8�#�b�9Z�6����V�I���0|{�ZfXj�� �ƀ��2���0��x�S��h+�-��A,�ҹ-�䌔���d�C�C���	��6�A�9�u|�0DL]q��:tYWZ���)x��U���)y4�B�1{�z�h����&���{"���|dV�^������'�`Xz�\�gO���^�û_�/f��U��Q�b��=+�N��6�p��>�#f���Gu�n_3,���T��:;#�M�Alhn0����Q#�����3�*/nIVMGo֧���)���y�L:А6Zb��
H�Pb
vZ4D:7Q��`��G&�0VKxIBF�]D b��ԙ���?R����MW���6�KO�Z�pЫJ=x[���m������)��D��G�DV9NTkK���Η�"�vN�ml� _ �a�%Ǽ��g�3�Ѱ��$��mi��)T3h]-tn�fC�0Q�	�\��VZ!���3�he�y��5ց2!��yȖF�xى��rC����;��9'��x�!�;H�&�¤r9� ��mw׳&i�k�Xh���a�&ʒ�b����8��	q��-ʎ��^�N4Eg���.}�����W��p,�'`q2�\Ol̓7�x�d�]{��S��y,5�G>/��Ȩ��(��j|��o�p$�sL]���B�v�Q:���Ŧ�d�I��s�]F
q�MN����<����d]��h�̏�C�4��ԝ�d�g�{"J0q[��QH؍h!�݄�'�;��;�|��|�Iۻ�TY2X�m�8@�v�m��Ɍ�%����H�}Sx+/)�T�
9�ǸX�y��#��	����΍|9A����ϚF������?%h�8h�ʒ�-��{'�� C��jQ/�~����O+{����Z�h�ѽ����!L$��y|�=P���ߵ~u�.Ǜ���d2�х�+SI,2�(�)�pGp����c�!s(�"<��]B��rԋ��q@�z�^_��3X�<p�Щ��#/5��0�%@��T�	W���'p+���ݎ���wI�ʁ��?�3��``�(���B�������mͤ�t��یbH�3V iڡ�wLGY�_(�T�۱/f����G�ҋ����&�>��9��-�Ǩ�i��&;�=�J��:��Vr��,������7��o�$6���N�-�e{W����`��*��*�e���&5�?S�:zBl����a�x`޶_˚ԹAJ���r�ap�38ſ���c���|ߩªV&UrJ9�}uy��w
whA���~ۆk��*LX�%���e����^��9B��ʧ���y���)u�������B<�6� w[��(%�+��֚�ǈY���(Bn*{H��oC����<�g0���B���;X���Ω�J�~(��x�d�(����^���Mo��)}��@�F�#+��q�?�
�+שX�T�7��&j��;�ʀ�����E�Ly�e�5�R ,-�tO[�i��ŖHeс)�L�����d��"�K����z����͚`ts��T�5�(�p� �|�n������'�����D��,o�"C�KG]�G�T��d�Ń��LڎAa���.%��k�ZP����!�N�ab���1H��%V�7C�$�Y0h�It��%�1�6h�z����9j����,��ے��mÌ@9���/�"�%ɣ�"?�Y1�$'V���n!.@G�5LK���|Fˮ�\���U�|��4=��J��\?�fJ��R�>��doZ �ԡ�W̱�*̇����9��pk,��TÌ��l��?��_?~!Z��ګ�0�4�T����B3��[	B�s�i1��}ϻg��iA�ޤ$�lw|��j����� ��l����#Vl�<�|UC�f�Y-3Z�e~@�HSH�Y[�J�8D�����|~�������w�.>�wPe�U(8Ң6�qai22�FD
\չu�9��pdD����\y�]��0�b��oya}��5�X�W"�qm`]�ݔd���NZ1�x��kp@��>���2m���U=�g���m�V��l�9����BE��� "�U:��v�qM���3��|)zy���F�u|)M�����m�X>�q����Aļv#-Ϲ.��)%^���׺����Y�Ҫ�,?ccP��kh0`��|y;���N~��c�f�'�G�UE���w�d�oJ�,3��"��G�^D �7a������K�*f�FQH�I�d��UP|r�&t<�� Ʋކ�:���;+�uL�������Q-��s�/���H1��8�'�'1Q������,V�Z�9���%u�mJ6ݞ�>�B�)��3E�*)���זB6�:՞0.a��+~��VKH��d�1��ƣ���P6u�IG�8R�Y鼼l9�,�r/�\��s�]�+
p4��ӝt�q+�BpG���g%0]�������0C��^�ʥ�+�X%ɱ��_�,+�T2P:/��6����n#��M�:$��=/�����	�?���{uk����F�b���Z���["нZL�tΰ+"����?�����9�K�%�,Ϳ��Z�i�Ə�aЁ�Y�)���%�u�Q�����=�=#
���:L���cK���|�0�����2������$j�S�O�44�JfA��<�]�r�uX���� a��>����k�}�M�����/Ry
e��[���m��j�F_y�1&i��剗Ҍ-w��^,p횎�?c���!�7%Z1f�l�,�=�[y���哄�ԎK(uW8�kW�Cy0]Xx��l��6x�