XlxV64EB    48bc    1290����>�̕ւ�����v�Ĩ��t��D�@֞PG��TC�m�ƍ1brAG1� ;7e�U����K�<��,E��'��(�)U=�P���%��=č�K�1�P����E���	vݚ�4�{٨�V�7>��C��fma�xF/��q�g�+j� �o��:*n��O����M:'��Wfl�'��thM�ڤ�؏/sw�����rm��J�D_Д!6$)m&�Ghq��ϣ
�a3?������Kˌi��`�VrgO�˸�{�u�H�~D��oA뢿"��9�0/)aX-g��t~1��..]&�1�tG5x�F��A���U�K�FKd�jKޣ_��~$l�����1� 8流�|��q:5cy�O_������r�iar#o��*���SP�����C��`
d����$���t�A&���i6Mm���vۯ��Yt�6� \:��Z�}���zJ�&�j��R;����nS��n���&�-�ό��K���->t��G��g�����䁏5�����=D�+�S�'���3��Eǭ�1r)B�,&�$� ����""gz'��vNY�;�E�,����v���{h���,�M�2��/'��;���~U�A��w~��o��#5s��f�@d�0=���&2x��Z�������o���!����ڴ�E潘�h��ڳ��5�coH�$��L�~�������Xo
?�%bZ�_3"9p��9�F
U��l�]`���rL;�/?W�:��H���V�[�0䟥�&�'Qݬ�r_��h��A>�:VY�?�<uF���w	МP#���Ț,�<[��O<aR2�}K۞H������$\Ag��5_�am�Аgd��I>E��������85�^���Ld��(��n��F)����1#�?l9�	X��
�u�خ�n��(�wm��Ȕ,եCF�Nk�w�Cc�Ρ���ӻ�M[�dVi�f��f����0�����I>N?h1���YNQ��GXD�#Mc�D��c�
n�P�o��QTJP�K/em�C�2U�}�}�O!2l R,e�q�0���������kL%yw�8:���2$��"5���B�W��Sf0&ʴ��) �'��&d��y�����</{-(;��Y������&H�Cm�ʣ��SU�����g�����-��_��a$�2�l4%�.�*�N������ )��� �b<ٸ�4�8ۻ�TB\Yo6�m��s�X�z�G(2��lQ�2��@�a���dKK�s��sOx��-RX�u;�D�b��3vb�ax�����/����v�W�@Z'q����p�\B>8&Ӆ^��'�)Y�A��\��*co7���*��=a�{a�(���3O�$��(�v�}���l"��JL`��zn��h�(���V7�O"@b�\J���"?~w��|	�J��{F��m�.���)�*d�H�.���vh�)<�Ŭ�z�^(�e3�����E7ާ>���cXBb�G����Z�i����kH�[i�}[cm�^�Ԟ�[Eu��}������{��0����ZӺ:��t���^zk M��"�Tӏ���ȽZxkED5Ђ�U����[� 3��[����b��+��C�P^~/��R�)���A5Gd�Ƣ��**� \)�*>�V���Tx[oQ�� ��;nW� �A2UTI
'��Ut�kb�t�,�v	MTοv�����;�0MT��Ĥ��)�?�R��'�!_޵���c���祅�~�PgӍr��8����l v���0�"�"'G�p̐ɵIf���
���eK"I�ݴ������l1�����<�Qd��D�s���h�W��2����h"ӆ��^ T�f?jpF63S�������I�Jm�g��=ץ;�0���2���w��c^I�v�� �5Go���U��k�VS�6f�f,q������������r��ۗh0;[��:���'PY��mL
�T82�X�0���2�����$�3h��p�-�9pւ���wM�g���DȎє|�KwDZϰčF>8I Q7+�+�;����o�@��{���G���)�v����P�Y�1{��R��b_��1z=��O�k#��<hK���¸cg`[KsKt���?m6�`��I�.Et�
r��R�/̣dR����u���L�u����q�$�f�dC�[Y��UkcScm�'⇫���qmc�u����;���.����xO��B`�u�b1���h��9�H�VAQ<���M�B�DC	�x}����ݻ�lڼ��}�K-@?:kZ_�H��a�eM�qC!{�[�e��a�F�U���T:I�λ"2�
���\�u�1���^���{>fvG$Oe�J7�F���F�W���Xbs)�9 �r�c��ѸAp�L�1�O ��3��>Y�� ���hY
L�F��5�pu��+��;�ҏ��ȸ�@	~���Yw+Y}������"��0?Z gqä����S�Fz&���~�s�gO��'� ���j%v `F����!9j>����]����Lfie,vA=��K+��2�w���	S�I&5x���R����STu���2����O���t�)۩4�+��޲ϼ*G!|ƴ�����"<�ve�Uɬ�2D$- �bHX�#^k{�U&R\��!�$D�d#W*c���Or�����$G���[� c1m������0E,�$��*�R��7X�����TJ{���x���������X�:�}Qf-�.y�^���
pb�vF��P�(۟�xJ��ft�z���a�sI���ޒ�>�E���\�-Ïů��K<�-U��И@e��O��c��z5���O��ȫg �y�ާ7?��G�[�{��_yg`��T�g���$u����O��;~������;x:H�lI���r�_d`ǳTX�!�-��P��H�i��p�������[�a�O�����D��)|fW�*2��X�]�e�Լ{���%����tA~��75�'�����Y��FQ�ՐZ!Y<D;H�ED�B '�4��mF�G����N	�TҦw�7��FF�����Ҹ�h�*-B�l�&��Z��I�w�YO��x�¡�VP�4H#�����6����3>��sE?����{} UU�$��1D����9]�k�� �Q�,N��� ��ˬ�==��F�O8��2��zl^zl�4�qxѯ�[l`,��T�E3����̗0<%KE{�V!a�r�۔��5#3'0�R�,G�o��8٭0�޴-[�k �p	$����F5EZeq`_ԝ�ق��~�E)�P���	,/�w�����(��G<4�;�9&r��n�&y_GW�yZ���A��a3����[Τ���s�̵k(�c�=�Z��ė�p�<b
@`O���趙C@�|��o��E �B �q��+�r�{Je����PV��G�v'{���u���>��N}~���vY�u�'��O;S�6UUg/m�0b��G���|կ����p��/I�a�(��t�do�L�Ś������N)[Wy%�B�����'�Jϛn� ��7|����UY��X�U������Q�Lz����Ҷ���`Ha&��!�x,���*�Gpj���G�	�S8Q<q�؀�׆��[��(K~$2��\~�3�^���)��5�]�ܗ��:��?��H{��B5}��3�e�肗���7	&��G����pk�gx����@���Cy�@" �\=���C?}n�7@��;y&�U%i8yT�C�!y�1ٌ��`f����y
#�3�5xI�O�:�!� !����I���D[ݝ�U���3�Z4��S}sP��>�5���u�gR��?I���Z��H�R����\X����m�
�a)P㕕MQv5���{l�:����zR��\�b����p���U�FI�ʲ-� �%��TV.;���A�qU}����"�wJܜl���["����P}��p`��!zՎ�	a$ـ�=]E��x��7��9�� S���fx=�R^�J,��:�u�֐|v8��Yy|�Ԁ Qh��jC��������lȥҺї�즟d���z	�Uuo-D�l�-1�N>@8D�GTh1e�Y�]�0H
�����ܽ���{i�yh-�Z��L�>��*�� A�Z�h��1֣���	�P��,ݧ@j��԰�#��XE�_'�a�/�
N	Ł��z�^��є�cB�4��i5��l���y�c����b>�Z���o'��zC9Q�p�H�D�����2@�W�C�U�G��l���2U"���q@���Hҁ][�@��O�>96}�h�u��s�@tf�;���x���-������^���`�*����]�������	�MKd��,^�7g�L�5f
����>���:���VI��YoK�ܠʣ��U���E^���D}U���>��N��#Wa���3a��������hP{h�Vų����7�o�3Y/S����O�!jb1
0F���
��N��k��m�^^?sS����&��k>y�����{L�.*T:o[��tM�H=�!{Bu{��������r�9���۳+�#yA<qBa˃���/|4,�I�Xl�����I����i*5�������8V>���T�HM6D���[�k�̔2�OJ�<Q!*UVRUg�qk�෡9�[!�S�5�b