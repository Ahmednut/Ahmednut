XlxV64EB    212f     ac0��k\1����}q!W7	H$�L�|I�����ox��XX�=�7�Rt`N�s��:Մ5&�����������,�y���䕻�|l��Tb�/�ڕ��X�gF�k�=9��​O�mRCff�Ա	~m7�w�,���[]��5��4�XK͒�F5��������w��W8mv���U��0�_�L7�HiTS�
kJ��Σ{��j�&��Cnp�{�����/­;��1	z^�rG�zC'Y��F�N7�9�J��x@�
a��c�|�wFG�Y��2�
�M嬾\�"��b�,,�����8
�w%Hc	�Q��j$�p�b� L������u��M4��� .,�	��(%�N�찲U^s�`��o�5v�cf-*��zR�\������r��e���$pJ==�z��mR<r�}��t(C�*�r:�G��i�Q���/��=��ܫV�'�ˬi&��.8j�KQ��ÂY[�A׾�;���p��GI��ec�ӗ�r��#�Ut�V���g��e��XR�$�0�^9��)���՛�%���O�yg�����q�Օ��*-� ��#8�h�$���X3�����MIDWh]�v@G��%��&a���9��떫ʃO�Ք9�t� �����Z��=�;j���bx���*]�6f���;�TY�������6Qߌ:�sR��ѳ+�{�b!٧m�}D��+�M�适a��=�̅�Ft��kO�/�{���d��Q����kE>|�A2v_��@П�G��/���)0��"+d��œ*�L�.�������-��D�~de��X-"4��JQ�)��@W��$��տZU{ؽ�r������P�-���v�圦��-\��2�`,�FG8m�x�&vǎ`���1g��M|p|���]��s �
�����L����3�ֿ��A�,��ۈ�f�n*��*�d�:͔����/[V�Q��#����!J��&��6M�L���x�-�b[��b������Bԉ��^贯�����l���y{'�&��v���@�~�,!!t�|���c�5%���O�i�4���T$G�[Mр�5T�}����ʵ��M�����X�.�=8�-�Ch���9��́�VP)Yf�i���d~b��
\��h���Ȅ�	� :b.��%)��2�[L��?4���˯C C
1���
7Q�&5������8�'/�(60�g���@m%md�����d�r3轭�?��|�RR�'b��+�	 ���0�Q"�"M)Z`�MHzvTp��1@�T�ס;,
�44�U���l`q;sz�QrYq��0�1>���yw�!�����d��X�u�HҺJ:� lMh��wDN���63]�HU����m4�u�z����}�u�e=cC��ѱ���ϺRr�g��=��9-���� �x4ñ���u!��IG�ɕ&�Z��B)C��AV�U��o��8Y�3U'X'����/�7tPs�Ġ��R�V]��  �:���7�y��<����?N�YO��e槩��%p��b^~�N%K�>b��Q����:��d�C�ݞ����0���
���#��0=:~����+V�S�!GA����� Q��S �nA�Y+�w�u����_n�,���K�>VdQ�,xVR?�]^�z�����S^��O�*�{b��k�$u*�t��������h��[�\g�<iZ�Fz��<�vxM��A0
��#���k���½��T&�h��
_�X��ꤲ!�����y� ܸ��ىe4��-0��p �."Ȩ����XF'wv���8���a�C9���[��~Ei��t�@���H��������G���}+�l�R��]�[�Z�A�@h�3���i�A~��%q�KMJi��Xi�1/hKT�Zc��4�����Ve�U�0���wH�񺞒a��k��mV��l?�}�䵔�5�N�f�!��:%eg�MJ�|����7��("DyJ���l�T2����2���i��`Ԓ��T��l/q�`\�bd��o���گ��<D=�؂�" ��V��ԾPE�U�����G<W\�66!&����W���Pi��y{g��1��ulx/W3 B��!�/\bar<}�h�N� �`�s��wMDHoM5buL)1�U���+������љ(&,�y����s�٩[KJ(a�hLO�P�����X-�E�@ldm�?��3�������ހ�y������$3��?Z�5�����?Z�-�0eՉ������hdv1��"��� :8}�Ԋ��·���,�v���'¿���E��֥1���x�s8�lJS>���H����
�=
6u��xJ�Y.��X�Q�9�{q�G��q��2�l�d�̹g ����e����C*5�Z�A��@K �ƃ�#��i��ɒ���uB9�+��ߔH5w
׺�����B�`y���Eܯ���/�E$* r��y�2�[���jz���X�?���t�`݁)bW^��S>(~h��i�u��f����)����)����*��U�}�ֻA�cD�@M�b��|8�0LZ���u�TZk9tLxr˘7ѷ����p���M�G)��.l���PO/}(M�����zL~�H�U<EK�$2}�wX�F�� �.]�����!P��F��E�-�%	-���OpHu��}�V�T��3>Sa�J���C�޹s@{���y��f
