XlxV64EB    fa00    2e10�d;�<��Y3j�r0�x��/�P��p~0��Z����P�jSO`�p���}��H����}�a�v�@�Fu�/H)H�@lN�!���H��eY툁u���;=�@��
��+����(@V�����>DW�M�	�d���֝��k:�VR1	b:��խ�#o�#��Ѫ�ۏr�^��$�{L[^�dp�:Bҍb������O;o����#�;����`��es(�_�h�SM�2K~��[�f�Ew������YĦ����A���ϼJ�,&6�/?;�տ>z���\&�C�*Ӥ� 5R�$���M�p��;��fV���s��1�+g&���<0�6�1����a?����6���G����5<�Z��@�� V\5I�_���@����Mg�����Ĩ\w�@�5
�@�/Kߛ��aq�9{&�?7�h�Vq�y�hȞ(�U��;�?�5�s�-�q��?�_�g���㴹&@W��5�����n�cs���<{�Q��_�����>�Z Bm(p����__�G�P&C#�y�O~��_�]�ќ_g����X	�Z�"�](�w���J�@ݐ$A��F=�@:�Q���!�'�c0�H�SŻ\p�˲����Q�����1��׽�`k��f�Gע�
���
��;��3����-����,�Ep��CB �.f�ϟ*�<�%�(�?�T��"ɋ�q2�a>�:�9V'u"��&<ͫX`9t��[����orA�����Zej�0�)>���>@_�|�
	�ߟ�O�6���<Cl:3MS�M�7����*�9����g��r�"~�� {�!��/�&���v�ɟr���*%����$Ơ�k	��0��j��d��u���b�bz����yZ�������wP8R���%,i�Ż���d���\(ش��5��f�܄B�Qq�U��"1h+3q���V�fnJR����i3g�F�ѵ���ytċ7���n@�Mc����D�{z70��b�Xet�K`t���_{�*$ ���!@�W�/& �Q9,~7�~��.D�JDS)���U>xh���R�JMY����LR,���"���e�G���@��1@WV�qv���=~$,�DF��F��\�	�+V���^�{)��H�׸�iE�\W�*����bv@��VB�Ш�ocw�e�T�
wP���/`��� ��sj���=��Oݵ��J{�M]��5�k��zD�ú�!�ƚ�!��lՑ��5�a�q��D1Q ��A�/.����L.�C-8j�.�Vg��-�r��8��X�Cϴ)�U_޼e��OR�MN7�Xq ���򣛵q�ry�k�Y�����ŭ�;�[Y�@�%c1*����<b��z�e�d����NT���~,�8�@.$.��e6c �u�ٻ2-'Ř����C\�*���P�V�0`�{�i�XT%
��w�(땫���;�w��>n9A1���OS�u*?ԫ�K3��R��&4>}���MP��o�)�I�`%o��U�P��{dD��؄Ϥ7�U&�v�9Wд�d^e�B��g �Z���Ε��n�h��E���;T�%";�(&f�ݘ��n��g]2�h���#��gӸ��cemы���(H�LV��p�=�z��
A5�5i�1�=B	5� ���������3�������ԩ��5L�@�|��L��D�H���\�w$rq�<�ESػ0��,wa9t2���{���Ң�p�2?�ۣ?ۘ��O50��K���;�TͶ
R��$�������l���b?|}�^�g
��4,�������_��:��jO���/\�[q��!�B(H��-`��_�ى7	�@̑�&x���	v
ph)�ps���n���ln�9�4+�G�$�-7�"��}'-,K ^�h�6P��ˋO��H�ue�!��!O��tEs�v�_U�jL}�����k�����u���ؐ��KfV��-���L23�����>��k&O�*�L����rE��p/���w��t��M')7�ݧ�4�����&�I�H�@�,Ć�~z�l�<�Ց8Put�zE��U�L��'��b)�{#m��lh��¯����2�Q`&Hg"���lqf����JT�f�dj���C-V��UV>��*GUX�H���v�=�t(�v���ben�R�&BE��mV/�b�_"f�2U����E�z,o��B����E�@o/p$b���y��j4EF{���v�t|�P]�����j#1��ݒ�&��(��cߓ�jM���k���2��`Z���d>�va�C��iҰ���б��n��6�E5S��紣�^�Ԃ�u�֙�nay�,�f7&<��3.�R����n���|yh �/�`����������x&p��a��NI~-�Xr�[���bwT�K_�!D��<|<����s����i��X"C?!w=�ɐ���>ˉؖ�D���B-��vt1R�UF{<Q���$�g�����]�!T�O�a`A�3`�������
H�*��F_p��l��'b�f9XZ~;�z����T�v�N#YP
P����Ӿ��\h#L�	'�5�@���[�"N��M�
T����5�[xm�NC}:V���c�<��+M.�������t��N�0�1�B�����'�,�_�jZY�H<V���t�t�0[`0�<Tf$R�M�#tk���!'L�4͘h-�PwR2d}��P���w�ܫB�`�nڣ7�e�qP��im[}Pn=ӵ�:#�O��1���NS���*�p:s  D��&C ��K��{�W�lu��ǧ�{�g�-RZ���B1��C���,aF����릡�����ʺ�J����-�&ЧѭQ??� �k]G �.��i�'��?;{~�Cf��d] 'Da7���l�� (�x�m��4�w|���q���V\��������ʇ�Hu!�	}�HXM<��-/sف��
��Z@yWo��8[�5鸟�I��̅��w��s^4f���0�aRQ����v�![l���vBl�L�����&^�7޹T��_��-� �{m�,w���)_i!����-��ffa��u{��m��TO���^z܉
}v���x���- ���l�J^�.�WG��y��i��U�q�E�% p��I��~�H��-0i��4�mS�LF���+Gqϕ��4��mh��lħ�=+�=�����xq6�}���M=�{��$���(=0��j\�Y�Qj��Ֆk?e�1��k�Fc��%6g��}�^m��W'�Q��
mS�b����\�*'y="�0��ԍ%�H&n���B/Yጇ��3㏓��\��'�š5$*|�A`l��0�*������I3,h�D%kT$$%h'}AzY���7���Fi�-ފ_�k�Qo�d�_j�T�ƨt�cJ�x�"��ǩj��P�.䑏r[*'��~�{-C�j�����3Ag~�ajzV��!�
M}�iL�����������VsZ����y�Ā�ۙk���+�Q�
vJu]�NG��L%S�.^���0Z�͸z��H�G��5!l��Ts�����7,5 p	���<�����~�
\����Ni�����2�f���+��a;�ʊ��c�ӓa'��Ԕ���=�*sVi�4C� RG�x�Ha�\�����
�����=��}%�A�{�t)%�zg�v	C��W�?��?e={��r�s�Fꉬ��t�W����y�'+�穦�һd����r�!���@�j�T+�>�49�(�+��pM�>���6Z�B7�sw��f���s�>��������(��"�<!�Jc�o3�|�o��&Ǥk�����%��Tx�O��[�P+tǄ�����W�S���%�P�'M��1�!W~Z:P��F�h4�U�M�+7KEGc-���F��Շ(+�V�=�j�&�G�S0�1�?ڧ	v��>���g>�}[ �I��v�5"�e���/3<����qν�;��A*���>����Ҳ����w@�(�h���0���]�=�Z�ODQ�2�a3�mTo�JyL���*1wJKk�&"ȩ������#��K~Ń�$�l� � "�\�Q�(8��X=E�۞����o�{����~Mm���<�P�,9���(h�JH�����Y��4�h�t�Z�о�������H��� ?3���)$��H��>s�;cy#�~��8����Sb7Y���Jq~X��`��ha�qKϝ��"�䃲�����S��W�v�ג7��À�z��㢐��_]~�d��h#�Џ䙕"��8.ȴ��α$���0OI|�3�9Fg�W�"����4�V�� >����]��
�L��D��t�᩵�%xV��K���4��|�ݻ4`�#�N��P-��8ӻY�H�uEtZ�@/$�}w�P�%�_���~�,G<�Cw/2�����[�m	j_zT�b&��[��T�z���_A�Z�3L�@��y�rA�/W�fa�����/|Pe`#��e��s�?�[�չ*�#�ac�U�WN�o����^���r��T��Ř���ے�ф�N{�!�C��6d�5�k�YH(��M�ɹJ�`�@�߬�����ө2I�7�~`B@�yò��v�V�E?{�;$d%��(rBK��.5�9�t�[��u%n�U;�l�~� ^e�q�ݓ�(+:�U�b�����T�#�*Z�J<JY�˞����_�ϓqV������dեS��'Ê��]g���+s�N�k[���N�M��[�f)���-R����Mo�=�U�$�[9��g��P-U�\����),4F\D�%�s)�lr�����!�-%h�>O`����l>	���8�7b[�(����D�+��A�l�����"��� ���d�Q�$�ﵗ=�Xx�5��>�g�����F5��0��K���o:]};�".���(�|�k6�������)��>����j����f��BY���G���T�V���D�?�j8�~��r�ò�q�8~}� ��q���42d�w��z�&�j˧�ߠ���J,?��23��D	y�qC~�+��EX���h�;(�G:Dչi���>��٘ƥ{}�:%�� ����u�%��{���S�3a��%#�޸.Z�j.����daD�p�.���8�6[��;A�d=�aɏ>�z��G;��^G� ܳf8&�5�F -h��Έ%x��:�����S�DJ�H0ݏL�,(�B��ө����U��\� ����-����>4[�]G`�ϙ�}��Eب��K��%�:���$�pKwipc|��a��=hb��sz(�dLYM�Z�7Ia����ؓe%��ʥ����@=ʀ������m�O)�3��*l��:�� ��Z�f,:0�+�N��Iw��	�����\���n������l>V�M�3V��f m_�2��M�S3g�~K��2ە�����
x/騗~%�y� ��^�S Л�5T��	Yh]�g�$Di��*:<�3��d���ؕ�7�sfΛp��-�|TG������q�K�X`K2�6��0����6nm�bNP���]�`;L0����9�Y�m��>t�5
@1��0h'�KL��oK ��;_}!-��]�����r�RpM��*7��Tx�@VR�+`s
zgp���>�w4)�\��[C�V�/ZS�O�CFnA؃���*�*�#���֮W?"�p<���y}���b^H�"u6:ؖ42=�	N�o�ӻ.�g�{�<O�E�np��'\/����5�
bD��Y�Mm���q�}�IY­����-�B�5�+��ֵ����q�jU]e|B�a�L�F�N�}��F�k��X��k\%D2N��������­�k��~�v��Zp(�[�������{1�����b^�zޱ�n���q�<�����/���^�x����@5�N����zqAF�,>,�q[�T�!��t>�qD�����_W����E6�~@�T`aL�-���/s�y@^^���� �m��N��r��
�2�/� �C��⻓��Ȥ�$7����b}E�{��0K:�p�摷;��Y4E�Ǻ���eZ�W��b�ػ�vO�>K�>Pz���(�BT3˕�Lom����PYeL�]��̥T�u�zN	���m�fk�8C{=t~r�(��
��#����
\4a@$���0h<I��h��
;^�Bb�=O��Ƽj�|f�x7�ND�H��_n�2�ci���Q�IzA}�t�b��J0��E0�O���.(��#��F�ths�_�<h��h]�4�,���қ�l{V,���.��5�p�m�'8`MzGQj�q	�u�ճ&r[��1�݌� / �
�Ϣ����@ij��H;i��~�K�6g�=������]�Z>�G�f5�.�$��o50O��i�	�.���R�Z�y�Hy�!$���R���]�(�|E\3g��+�ͯ���D����]��H���3�7$�(�����fk�JPu���v8{��*����Ц���)�u.�tt,B���D����/C �%��`L�fdu�����;���Xx:��g��h�����AJ�j��l��<�>A�vv�,�&��7+�f���G�4�����n���0��܃�8�K|O��u��v��t̶^3��v˸N/����^
��Җ/ Ͷ����L�_�6q2��C����b����ɇ3���+�!�<R���|�Y&�^b��쵗�6�0�μp^��{����L���5n��]�%M>��o?�}B���rZ�eI�Vn�}b�I�Y*�4ߎY�%�`X���<h)��,��[\�u(s.5ma_$�c%9��_L�Zf�Y���W��H�!u/�{��t����PVVȋTL�}���������������ӵ�Kkb��e��7�V���X�Z�>�a�F8��Qjȣ����CB:��pPp��9vۼ7�;#|D�/��5��4ܬ�*�⇽�{�,��k���^*��i��%��C:;��g�S{�y��c�L�A	Z�Z���]��=jiQ�]d�B����G:����cA�qo�Ҡ)��ԧ�7ËO%�bVp��J-�ƞ&]e�	+�W�+}(�WR��& rt�W����?�e~$tw� G��0�{� �T=>���OM��'V��%��pv.�"��Z#�'�S�yPt�b�ܡ�_3k�=�sV@��t%��2s]�n��-�Wx�zš_*�MiB ��6=>yZ
M���MK�ĪJ������TV�$IַQ����eˣk|8����[~mF�u�(�o��(�i�d|���R��qL�Z�� ����g+���N	��O�o8rt͉��]�C�Ay<Gs��Bq�:������j�܅뿞{��!�tC�L�	��L�v"�Z3�z�I[����t"5
�F�r�b{"�����=����̱�c�h�z�G�8��ʗ��:�qY��_�"�Rk����P������\�BhF�'�/��
o�7q�|n���qcq�����]�������,]��� >���b����7����❴�������/75�	V¼�"$�G�t�&�蔛eoKU�E>�B��8y⎏=�M9{1��,����?za�^�V9Zg�"�!2눒��>���I&ke?a�D�^	 C	&Z��6ܶJ�j�dl�����HK7=���B)�'K���jtM?�n��V'������2��B�ї���_�=��ϵ\	I����:�բ�$\���#/f���f+^J1����Q����/'�����z�B��.���mՉ�=U��LӰ�[����Ƃ�(D�OS���_���k��Du�o�n7B�.�LW��[n"��k�ck�w���cOd� �닱�~��iÎ��!��m�h_XZY��)A��J���9���(+޲P]�O��r��3��������J��nW�#�G0�
�V�2�#[��A!�E�i�ʷU�3xw�iw`� �(GǊR�e�x!�+��/��]oK>�MŪd�Bh��3�^9�{>4#$Ƽ�q�c� NAw�}���dpNջ/���	ŃF�?���Kw)�0��޲%�.���v�\v`w@�T�-�������qs��
����_���vv��[\��JӔ��:qR�B��<� �K�3��+ ������/c�*�!�ώ�,���K� ���cr*Ӌ�5zׂ��m�RϤF���@)�j���U��n��~u�{���!l!^_�tI2m�[�%?}���su��19필xP�4����;u�?v������Zyë��r�W�E�����4�y0Z�����6�е�Yܸ��a�4#�G_-��S�y��w=(������+���S�1����2/3
iϛST޽(v*YA"5!�I��(I	�<�{���J;-�0=��s��f�B�(�����(e6"~��R�2�fv*�U���㍔�7���PԿ��QR��'� �s�7��,di������`V�\_C۰�`�<ۆ�Ǌ�T��F�ةye�#�D2�����Y���;���~L��Jd����
}�<o�"Kgǻm*/���ߥ�2��P����&ǺM�l�ۧ�#	g���ZTHG|YéA{S��V�Q髆O���B��!�o�o[	8��@Rͷ�(�QG�Ʌ`byS�W�� ��r�q�nt(8�H���ϰ��Q�ءT� ԡ碣� d�,+�Fy(/�<�xz�.d�=�Kma���cK�[}^���^�$�p�ȃm��`Xh�/��E	��i����(w�V���@ �tNM!�x��]��_c��1�,�S@SN^�\�b�a�.��Q(�6g��x���@�M�k����jy���~x�sR?3��a�����F���ĳ%u��a��������9Eǿ�Ӕ��������;uq_��#K�xzN=�v�{^�˘��r�2%�޾|5+��Er�B$��8�Wu_���B�U]��)^/iv*�2���Zp|7�`ғ�($z�O��H�9D��?���Y�/|�]����w	t����H�p�P�N�����5&%f7}`*�[Iaұ���dG�rmKoA��z8��efx82ٙ,X�|0,�k�*�]��t��B@9��"�G�㻈	N�T@�#�
�K���a a��!��Z�z�������ET��	)1ݘa���\W�X#7���M*�5�#I�w��̅�2�"�r}8����2��Ɛ�E�i�P��l�"oU@��q]VL�Sc�G5�N�-�'�wA�<h��h�-埙E;i)�:%�rc������Q�O���;�Y���[��ޣ��І1uh��1�?�U[[�'�頚S�c�;JJ�SZL��S����~��T8�
�`eyP�j-�Db���Ճ^.�ʳUV�3�Zk�$~�=�
�zw*��pQ�HIq�b�����p��Mۯ���]>�Z�`۫#i!h��]��+�b�Em���ZG��#�:�Hû��d|���=�rxMȾ|�E�;�GhK��O֢���,L����qg)u���z`C���m�s�� 1�80������֤��]�\u�3PK�L
���ܔS�}1���O5�ll���µ6�a�n��hͳ���1#I}�K)�6$���>{�=�Ǭ��[f���|������P�s1-@�o��Kmo	���>�v�gݧF�?�.V)�1X(��k�o�HD�ʕ���fbS�3�Њ��!�V�R㿿����_j��:X	+��:������R��"�(ba������NM�_�Y�V��D{~덛]����t���J]n��x�T���|u�>Jx�8������:�~ͨ7,��N\����ӐǈL����zS���'R���Hd�W���`z�$�\A	�(I�0^� ��2B/��;���JNGV�F�"�wJ�4���9��V�Oՠ�4��:T���f�E�7�v�'�Ɛ��zՈ2�D(���E����O�J�N}��4G�� F��f\��#V�hͷu՛��Vf�o	���4)�@�t�S�� VR�/fUX�_��:jM���s����ᵭ�x��N{X�#G&3X�a�z��&Լ�o���T|q1Ό[��7��,�%T�.���C�{rZ��=�r�)r��m� X^|��z��詹[b�Rѣ!�^Q�����[����3-�� �O��#��_�&3*+xq|���d밠��h,��5j��;�8���_dE�ɑ�ے��w��HWvd��p��jKB6Ϛbf6�H��J�eT�c���C$��+\���3~�9�x�Tه���D����\�
Q ޙ�w.Ȋ+�ʇ4%$p7��
;�=`��5mD:�T�=�\�4��^(+"�,�^^9ɔ���M>{#x�L��M"�$:�����*�GY�;����a�Vu��,=��0�!��-�N��`1���+�� ��6&S��2	&�@�O[�M���2�ф��(�33n_d���P���͝
'�56Pz�N��H�=*?�f`���.��J��n�r�y�,��#ķ�	�����'�a�U����A�����td�X�3UB�Sj��Kw�ǯr�^ѳ�M��3qO "sa낓��N3�N>�8t�� ��΍�YC�L�(n��t��a`u%��|��A>�t�R���y�����庲��+]FB w�G>�rPXY��������f��^4��^����O��Q��](�qU�g�^.���.3=-�"�_�c/�4�@���^ŗ�����B�
���z�w��q�{�s�G1�����"9�ې6I]f�t�6���c��Ll�m�c&I
2�����}|�2U)p��J��󲓷��x�#OJ��T��<%�ߖ�����T]�L?C*F�p)����h<``cˍ��q١"���!���f4x���NI�;��J�{�<��q��K%h�t�ei�*G�\ֻ�c�C!r1��վ��	P3
e`���.?�I`1��m]����:�����\�Z�tw���h�b �
F*,�H�R��ɬ��kkw�eT��["k@��M�\[�W1#�����mm��x���ºQ}�Z�̥��(�������9�X�5��97����(�l�y��P���@�A���m��[_��������qa�����{�(�h���Y�`<�LD)��ΉZ��h鲐���>u��5� �"�*1��f<S���	�dZD�|/l�[E1w�ly�N���Iy�`DJ�ѥ���.0�l������5�d�AA�s,����X���ve�pS��H��E�n��� ���~�8Q��<D��	���R���ż
�ղ��"�s�Q	=�W;�	��ӊ��w�%�G ���5�K���w���H�����0�����x~Bb=Ь����6?N�$�j
=��I(��B�����m&Y!֑�f�]^=wc�ް}~`zB���^x}��έ^�UAF�zi$���O�i�z��_Ys!NpV��g���p����u�|mJ�\��,Ja�0ة�5��,�B3E���!��gth�Gv�J]iK�:r�HeD�T�ۢ�����؏	��7�c)�ԼG:#�{�)�᪲�A��o�i�{.��1E��2��Q^oO©ɫ���1�����u�mH���*����z>����~�By��'�P\[���/!q��9f�U�XlxV64EB    b567    1ba0�Tsm������cv.*j��b�����Å[�|���5[ek��/ H�4��M7�'��l�?g��uO�7��Q�&� �=y�Wrf�͢S";��y��f�ß�ؘ��	�Q]\��Ha#�p��;�2L"� �5���3��A㓃Bo]
=, ��n/)%%&��]����quR��żlj��U��yеDU��	'������Jl�T�V#��<�Y�L3fH<e w�W�x\�|���������<�%|����珢�]�,�6���t���;l��u�A2�72\�5��yA�>�W�����
W9��}��H� ��-@U�ή	f7�w��˺o�¤������j @�2��3A�s3A1%����"f!E�2V��i�cvHֹ��?����cC��O��9Ef{-EOFۯ��63<WޜM!3�K��{�A7�*/�j4/���5�K8�sx�2"(�'��܍	�(4��
62�jK��9�������N�E��1�J���z���V���_�'P���f�hfT8�>H|0^w��D�����Y�� �ض��r$)��7tk��dU�>3��������'u h�F�!�!�9mb�:������?@WP�� 6_ۍ���u��K��m.)'�/=ܟ��]왌z��5�h���R�2G��jdl�����/+v]�\��,t����Q�x��W�+%Y���Zf�(=w����l(a.��Ii�x�!���W��-� �3; J��H�Zx���S�&���=j�Z*4�������lT#�ʮ0��ꌴ��B�1LA�b{fI2�(��`�^E*f�K��PHyN�Z�O�p�Jn��!�@�H?d(�
,~Q`o�E3��n����o�ĺ��z�� ���ČM{Tv@���W�v3��qӻ��e����RJ]��=�ܹ�k!�x���H��-���7�;������*!��l��Ɇ���͌epD�+c��*h��7��o}�>��e
�ѿߤ�;�������M��}1���m�����@������D���$�����@j,�"�68�P�k	��R2�%x�!�
��n���hA��V^g�T��v�o�:}O��/t	�s�u�@��[ᆉ6�5w�9�����ҏ�,��b��bM��Më?q�b���Zj�r	�۱\{N!��� �ԗM�o�]����Zw�:���a��=
�RZT����Q�bioă�]�#hG�f�K�p�Q��'�C�ɲ�m׬�$�������ng��5���6$�2L4��½����D�*��*9�ӕ��8���n�)h�[x�$�n��JV��t����ktq��#_�:D-��¡Yd �`6��C<ov@FT��u�$�5��)n�t'J6��^ ���h�&�1���|��q�{�E�%���]����$\����h�1�&=�>���l�zI�1�V��P���@س��1�G�Q�=�ʰ�� 	k��ɧ�=s�D��PƤ1�g����K�k�Nw b�dt�NF&�\�`�k@eD�u��O�y��U�j�n<N4cӋ��au ��] neE� O�k!)l�����o�����t����@rB�8��}(C���A��XWwڜ!�Ҥ*��U I�����4�<RHkj��r����s��4Ou��^��)�q����A���O��(�:G� 1�W�זV�KHm���hY]��_�zub�L������&�Q�H�M���䄬�S�{��������%<��f+���2��-1��g�A�Oӿ$G1�c�/'��_i�i�E΀W�:��|�l�!�E=mN���/>i�����8a�����z>�X���mQkB�����5�ٰ����ҡ��K�ouM��|R?�=����#�	�yD�K���8�	ӀF�lb��R�L�tT�
�gF�<{��+���z�G�*X_Gf���E��}�5�zHMdw Eq]��=K��nxM�
@��՟%��f�vMe`S�i�@k]�=Em��6�WCw/�-e^ra�}�=�>\#P=��ʹ�/���Dv�r#�����CJibû��p�?Ud����fi�J{=V�\C�`x C�,?̳̾���:����^�	ZQ1i���R|1ۈ/ˡ*�2�C���~��^����D����>�8�P�W�r32H&g�<�&��ǃTI�`�COy����m� q.�~9�p��M�'�Zs�	��^&��	��ԯ�3l�%~p���72�����L�[WջcVhc�(ل���I�F��(*�'���Pޥ��dgf���2�f�=��RB;��̈́c�p�8�w�8����qed���,@V�LQ��?O�V1���=���R9��ĩCʆ̸$Ë��U�Z��U�d�Y��ኗ�;;��#�N��e��
+*��6�gRT�'�F5t�۳�vGnby���C�� ��X�ЌqA!����z2)�4dxN����=ˡђ���Ȍ��-q.���׉��i��B�b�7~Rw{-�����sI/�.��77��n�Ysw�g���sc�אVa�v��_>�a1.T�rvnT���^��3h�y̑��ϭ)|	�J���"�r��oz��b.M'S	AD��M�X�cO!^~),�4~B���� �~���*��4	�>�O�\�]��I箱���&r>�����9$k�P�%I*��I��V7C��{�9�d}j🭢����N���{���"��;E��S7�q���}H)��Vdf0.o3�ט�F�|DW̽����8��mf�������mѺнg��Rv"f��et5.���U1�9��C��|�p�w��Xn�-x�'t|��z�)s�Y�L��</��N�.�_}�6��b-�V��4/ ����}�#7e<�K�g��v>�u٤� �1����W����y�(�8� 4�����`Us�V�ʳ�\�m��]6�)��v��a�kӗ��h����8��&{�m	����B%�e�xy4j�S�T���M�$Mb�ZO�́�g�>�3|��[���9��;�.ؗYf��q�����J�k�E����?�V��9�Gخ�ЎfXHD뜵��sS���3����+?���al�>�N�n�6�<�L$wRO�#��ξo��T�z�}N��:c�&�I��d�Lv���+î�s]>f�}ꦁ����B�t}�ŵ�7��_�ݿ@�S�dv��
|DBb()-[A@;���u�ت�6'�TZ��������C��ITd!L��[hɳw}3l�ȫ�ŦJP��nv�>�,IX�QZ�Az���-v��QaK4�Bz�>1D��}z���Ղ�bK�4����-D���\�������z`�~�X�t�/R�dϨ�.�ŭp�Bh���$A��31���!%J����ͯ���}Z�n����lbD� d	Nu�r(quE��h�:�朴Gd�r�h,��Ί�6��7)��3@�� ��>�{��@��`Rr�ˣ�B���8��!�}J���K������y�^���]j=-ۗNߛ�=^�AA�v�L�t�q�pB��pT�6�^�쀤��BC�RZeݞ!~�SK�ޓ%_�|�Һ�{���� �3?�ӄ�3~�Fd���-�53� �Ƹ^��SVrR?�a��WI޺��f,C�4�r�R�{� x�7h$(��ơ�</�?�~��UK��nŃ;w��G���(Ĳi��"R3�^
g��J%t��UH��3���� ����Ҝ@��D��OF��QVn9{%\�%����8�x&�~/%��A�������>Xa��*���t7��i����}�?�p�ȴT����5w�����{)s��(3V��K�	#q=N��I%:6��$.*���#ڂmqk���	Cq�k����\p�iHVKV�_���mHk�h*pTc���4�&#�1D��!�jX�bV������Ā��wh3Ww�3���1�,-�C���gve�#�� J�$!(Y(_h�k+S2��
غ�]�"���������J[��^��̳���s_��ZW[avFvV�J8gO�'>�= ��HSAIK�jO�lQ��J3��ja�7�E���v�_:Q����A���&���vHAP�s��������6��{quwb��6\��_�ҬV]��z��t8?h5��`ii�uB��ۈ����&i�!�qዬu��U7�D�9)	)J��?4MB�\���)3���rY�k%�Ì�cU�+a���v�}����~l6acw����l�c�~�5>0=����i�v�����c]����T�k��� .� ���x͋[�����R�m*&�C�
�sQ}ײ\߾�
ʼ؞C��jV�"#��@�M�|����c� �<����w*��.
��`n�Ae�E��hM��A�!�Y��Xd�����0n�Q$zV�t����%��mtk5�0������cp{{~v�}j^��K��^@��r�C�\�	��q�iZ$�vX��T졫 j��y\~h�H�*�̃9R���C�X����56���>���d`�v�L���d��F����PBȅl ����	!�+m�2Wʹ�R���) ��X��BX҇K �.�rs$h���h`@���g���H��Z�XU���D�@1b�Ӹ~�#"��AН���\� Z�g[��8*z�4��
���X��k�7�o�v'�	Y���@4�)R��l�{��3:����g�����Uy*�����ݢ��6��n�:�2�T��^����m�r�A>Rh4lRj���[� ���ԭN4Q�ښ?5��*j.k�K��8�`t���a��θа�ě�(�-M�kȴ�y[�%�0$��M��po���f���%�fn"HI	W�]e��~��Ћ�<�9�ҷ�+��(=K]���qʲ�BU߲��s6x�!|������������@�	#-�O�Qy�m���ؔ�}�+��;/0����GB?%� �i�:�|����l�]MC��Z:s�"��O�:^/b�;�	vX�O�G��fd������LM}H��J�"����.ĝ�ͻ�A���F!�j��B����J�(��,.��+C N�7�GO%&T��p�Z�ݘxA,0\��@TE��'�R�_Gs�ZI�yy���=��J�	w�w�n��ք�qI Ue���@�/�j��e�z�/�S����0i��B�;�H�^���<����*o@����e����W3�qO:�o�ap�����>���H?Pj3�4U�Br��P�g�Ր��W����Ħ��ӂlU#H;��7��EĂ�H޶'���.�|��dm�G2��� �!��b!M\�����/��M��?��(�0�9��&�R8�I��S����Е,b��<G�=����W\�ڰ�v�����i����C�D^�NoO1��,�n�W�X^���@!�w[�����9�]07�	��Lpސj��#i�����7�ퟄ�'=�_��r�c�0����A�f%�D��SȻEHEj[�C���Ɵ�H~�!��q�lZ��=[(��ً�]�8���l�����{~8pTh��:��w0�5�z��u�k5+6�4�
NU����3��I��r#��+S�p�~���ek��[��Ʃ?M�Ϭ�h��2.���\�f+qk��Wk<<I��K�0�VS;��4|������r��ge�3ƕ�5In�BTs�,�պ��y��X�3(�pbT������l��)���V(e�G�q�N��[8����,�{Lth�
]Y�J�A���c4ۋw�'�Kmm��r��dȥ܉v�<���4z��:w��0h��~O�O�`��F$C���"g�����C&yK���l9�l���
�q�QĴ��k&��`�>�V?�3�'Ӧ��#� ��?��X_�U�x�ă�R��(P����}{A�?���r'��F��*��`��E��	��xr�0�I(p��-��Ͽ�/�k0�ԉwaq�0���#*ET#+�p�-Ǽv��Z�0\�'�����廤���Г�VB�a���Kl���>���и3瀮����}߸C��.��s��)�r�����_(�5	M���/��
�qr�/0���D�f�H����&S��վ�B^�A��<���Zʂ�Q�t��҆4s�&I��I[DӨ���=���IO~��v1$���yu'
�J�;�o�\�W��&�����S�i��ؚ��A�@4�k�mI�m�-��~���n')�g�MQ�%��؎�J�h9��{W!� 
��=���*��a+�x{D. Sꕵ�ܐ_�ZTE�i�A�RkH��<��K�"�'_�a���AL�{bԕ�I���p���&i�il�g��ܼ��Ĩ&oz_������T�7׶<,p;���x4�dJ��ۆ]�O�9s�]2n�S�w��K[�]�=����Mx�[�dU>H��'͈@qrĘςPҠ]͂��j��.^��a�v۰)W��w��a�&�����I�b
���
�_�8A�^.4r����媮
^�1l* j8^�g���S�Z�b��?&soK�~��<%����^�6\&����E
��qm�F�����r���O��U��B�X�X?����+at�z��A���*��E
97wݙef�.���Ŕ rS��+	MF�IK�  ܳG_����-��qa9���3�%�?�R'��5�Ǘr��ˇ8l:�Y��|�W"��+#�QW���ڼ�7��	���Ȱ�1���l<H�Ţ�m���o#�{�Lᆵ @l�A�3�L����ja�2r9FP�>}��UbP!�Ԑ{���_���uݜʕn~�d6M�j0��v7�!7hT����E(å�D�l��������l��j@�`&=�(�lP�Ν���"��SGL���eٴ�h�t��i��l* �5I:�� <��jY�$6�`<����+%