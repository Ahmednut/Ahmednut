XlxV64EB    55c4    13b0l�s�2f_��l�_������e�^�	IbS�b�C7TsK�4��F�ہ �hĂ0��?(�:����1�u�&�VD��l�ڝ�H�@͘��Z�w�~���x���e���Av�ƺɓ��C��(�����S5
�|�y曻�,�6�:�B�
�T��k)q��!r|6�>�P�˰Vj���	�QAw6ј����G�g��2Jߩ������l�y��į��k�74}�F�)���Ѽe����Γ�|�Q���)��TڰB�~�w�Κ����I��ܣK5��"�4�Cy��Y�>F(���C�����w@e����ɢ0<��6PO`�y��0ke�9�"���!U7��K��I>��w0T�6������c-��T*�щ��ں4DF �8k�<�҇��ұ[FO+�5�	D� ôs\��Y$��^��1MR��>�(}X�7Y���S�@�Em�-�#u45�����Q`5�U�j3b/��2������Ұ#�ҹ�9v��$�G���:��0]�I�)"g��DF�:=.�����N�NLn��u���ӣ	뿢�4n�V~ _(ו���]a���VW�.S�MG�n2X}h2�1���֋���֘�c�	8#C{�~4��>:ǥC@�J@p�7�$6l}K[S^U�i��;~>���a#m>�l����k�e��䮿�c��WL �8��8���{�R�����t�����+]��	0�O���j��h-��z�g���o�hz�@�?[��n��#���)��]�����T��7�Gp�9m�^�g[+�6�a.��Qr#��WZ����`L'+���v��8f$��h��s"Z�l�U���h���}g_��3�j���y��x#9 ��M��q�kӄ����u�`1�1�c5�%Q��<{��C|K���+̸�K���=牔�]up����JNS�i �H�2T����Q� �3Cɥ�Vo[%�[	]�^���cIo_�Fe�q^���bU��A"I���	���R����_Y��7N��}k�����&��T�
b޼E���^�]�H*��Qj�����$�x�&�F��#ȁD��{�&�5����r��"mz)�^F K���~>�����l� ���l8eTP����1v�	��:A��Tʥ��b���ʞ�-�!Y댾f����U�p��Ҿd���Mv�8{���P����J �Q"�g ��Sh�<�	��o���@<r��,>{p��^`���.4W'nnUz���[��x�"E9zPY��~�
�������㫧~��]h8C{c���Z��8�#*5n�F�U��G�(��}=Z�~�1y>��]������޿E����� ^8����*��+��f�K#��Ү���̐��
��st���Pr�D�o�����nzk��-�y.:ƕ|R{���[���KF���������x�}�q��?RƼhRZ��Udځ�5�Jq8Q���kX���*e�S��k5�cu�!d�����Y���Y������<ٟ��ط��|��R0O��$@ڻ�{ �̈́�ƴ5h]<��C�fr#��Z&Z��T�)��O��7�,	Z��۠ؗ~H�J�dF�8����~�L�24Л4Ā~X��_��W��A����)qe����T�π ���J��ޘ���u-�-�8�ЄF�3&_(�|"���^o�J'Y 9�.���+�aJ�Z�<���c�O�m;d�sY�4�	��� U~Ҡ;��Ra�+b\Y�te,�����4�^���%\��,���W2�>F� ��d~����/<�!�w�\9��qY�𘸗����漐k��JV]D�':�F�$n�f��-����gvhe��O�sC�S��"���+/<�x��h�.�n�ڙn� �4��m0M���L��{D��3fZ:�2B�cI�P���胛�o|�0��h�%z��1�R>��l]��Lih�J;?5/u��惖�Wh�h����Yr�� �꿈����>�t�zxbYU�P]��N���s���82k���/��Y�\��ѿ��1<Hyەޟ��'3|t���X����t��$'wxRc��� \\L0)T$��]^�o��F�3� ��+�{3Q�jK�?���҂:��y��6��H.���g�qB73�6f�.�2<1m�]��͓#+p��cA��t�w6C�w��lm��}�
�&�����gX�X�w��$�f����r\,]��Ij�~�A,��V�PѽcöteEQ��ꓚ����4�4!_GD�ؖ��~�ga�%b6������A�y�<F��(1s&װ��?J�?�_�K@��B�}�n����&�P$a1�+�?T�{�L��+2�1�خ�$�@"pTS%F����{PRA+~�Դ��}�
9HNdj�%��'�����3�?�Q�� �iܮ��5Ls����HܨȒ8{����?N�~�������%�S���ur�|k�/8�7��U�7]t���R�dG�^�"�v��핷O��56��B!ppMѢ>~��0UՈ��Pa�M @�����8AЙ�l-��;�sђZ�a1��5��R�^��9�b>Z���I��rW�}��EJ�DF���بV�����V���i�'�6�?��0=�����57�I}J�I�Yƫ�׬�1*����1W󻎽���	��'��y��t�.1��u�\�R���,�˃�:��Nb��$���h�k���Z q\RS��`�� ����� ���igW�ղ]eSo.(!E�fgwU)U3��M�|��A��{�,ը7c
ɪcj��
Z��^��=�Mg_J�M [! [�%�8�cH̴v\���Q~:���n�F	ؗ3�(SADQD�a3h�S�L�qۄ�P�<�����=�yARD���2lwC����w�`D��B����������ҽj�t  �l��8_ى8��8���ӒEH�tƊ��!����z������[+M�a��c�)���1��3��[\Ccʛ�u�zS�s= v�~��ԙa���&�<��+<��aC-�utO��b�rb���8�҄k2Z+o��qd�8�����d'g�c�+Kx��2�����as�b��a{��|��[�M�u�oz�Ͱ���\M�iӻ*����T/�Йv�<�)$(�(�� �3����%S��b�\z��+�����>:�"6m�yi������k�-!��@�ɟ*|�
��G�5��D{D|���v�47����w3����}�A���L�W�H�!������D̐�doR��&���U��E�8���F'�����*��L��B:�uóZ���{�l����%O	�#�����){�p�X��@I]��������qB���%2��q_@�1��_�0�ĕ�a5^ko�D�Ȩ�.]�ȿ^��mK�џM k�ӈ�WɎ��%�~Ln�����;�^���wX�1�%���J��(<jTQ�a/����`�:48<���[~/���!;z~q���Ad8t
�-kOg������r�.!��J����*N����k�u���E���	=�o�KFB��=���ڏo�y�HaH���¼�'�{ӳ~[IM� 4��ɛ����/�O��d�rE.��Khv��s�� ���i�O�^�xw�`����-1�;y ^�i�07����dg���+C ��A&�*��p�k�h)H;V�7��úZ���g���Ȓ�P�Ie��DU-�h��_��O42U�b��g)�(�ɐ�����U{���5i�yϩu�ii�{���,���R˸����ul������N�^a�y�P�"���wX�O�"��
n xj8�Lz�� ű�)*���*N+-�;A�b���
D0�^���[Q ��I��6�p���\M# ���O� ��F��^q��y��g��}%(g���VY��@�}�|���5�b(wl�:NP�:��'�k	M�'�d-_G�׻H!S�<�w�&-8��m��H���E��Q��ji�b0�E�����54��ɏ��;��B*��S�w��Y�7��ޚ��q�p�>�K��yVv�>Y��D�&&�j�ͨ���V��N_xo�'�S��&ot�c"=�+�K�����:p���ά��0�g)KV�r����G11FF']f���kJ���=��fN�� �~�4��¿h��,Ow�:8C��*kP��TFI�CV�H"�gw���S$@��(#�0������]�vf��yc�L	;��kVO���Gn�z�B䅥� Y'L�m\��Ǟ+���30�LM�'ĳR ��ϧ�^-�?�; 7�&�k�$1i�{��hϺ���=&fF#̉u����%�����6ȯ:�Q���S�ZN#�8�I�_�1	aB��S+�NB����,vo���1����A�4}��\J�ں���z=,�Zk�1��U��$�,���3��O�D-3�M�:�sF:_���L\[����!���V���<cfDR1�����/&���:.?��\����G�B:a����D�J�]��U������PU���Nm���x{f��@;�5��/�0O,�_X����FX��83��B4�N�E\C��#2����A��
��;e\%/�e�_�?�k��x�\�R�+Fڅ�0d���� I��U�6�'�ȷ���\�LƔ�mϜ��J�"�♉�>�@H����!޽�h���kw�fc���*�gէ�K����_����Z�n��
wLB�P_\��%���{�3�=F���C���E���r��sd�l��+�u�w�����F�8ߔ���.��u'%+�|�J��| Y�ќ'�.
Q���~����02�x����@F����4�,�*�^x�	�
�1���*�Oݢ��\R^}4~ЁR7�ET�} ����4����uur�=3_�Ow+��s���7k4-UX���W�