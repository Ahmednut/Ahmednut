XlxV64EB    239c     b30��l�%g�������?r�#F]{c��Q��Uh��wU��8�9��|��M������A`W��ɤA7����r�ji�u�c�x���|Rx��P�bV�p4�׊jp��������~�l����+^��}���cF�V�}K��̢�s�,�u��0R�u��銨�W t�b�J��"/��J?iF�;vO�����g���9����چN%^YE�O���#թF��r�/sh�l��Ë���mP�����i=����9��
I��''�S��F.$$)	[�2�Cjg�HZ|����as�k="����$�w�c��	:y#���W�����a��lZ��u���A�Mx�-n�9�\Q'S�Lqp��I��zv�<>qKh��{���m�h���T�,g�H��1h#9�d�c&"}�����5h>-
V��+�����U�<�1�O�(k�=��-G���nz�����/�vrm���5��C��wc_b���F����u�&����,��C�C@�3�ERC¸����Gg���~jb�TT�.\�.�+�b':4��^��ی�v����a��r1ݨJU\��?Eo���6����eE�4yA�1�h��ӿѺ�*�Q3�Kfެ��K0���bF�H��4�����J2ي����S��<n�!�gt� z�]�ϣI��@�b�-9�K�֐o�޼1�|g�^�ޅ7���ex���g�	$4}�x�:�e�4���`nHwȷ��!�JZ��xT�p`Qv��ؾ�6FpW���>��nL+���-ȡo\i���!����i��1�@�M|t�+�C�eK�Ѩ7yw���BZ�h��������
42')��N�$~�K���ϣ8F�զ2���U�SnxF�-�)���F�|'�)�%���6p��C��E�`;S�<#N��O�N+D�C;o|^���T�*`S>sK��!�NRð�~,�������������vMm���
X����\/;�AL���j/:����Ue�u�P��Z�}���L� x��/��x}�c��P�������`�jkATpmw@��LA�+Q0�&��<Q)9h��Lg�@��-��G-ɲl�)�>����m;��̾���h����������;�믑�h�&_ĜaR@u҆��`'��K�_x�+r lT�m1
���+�.���Mp�|\���	N�7,�|����[��T6�.yD�ʗ8-6r,��>|�@n%\:��Y��a�F�t����6�yy=���=n����{#��P=
xF�+w����{�#�Wf��0So�)�%j��dKqD�ū&��_�'\�9^ݤ�� ��r�S-�3�!�J�Q�M���<(e]Kޢ����U�v�ܵF���Bg'IHgRqV���ˡ@n��y�k���Uᤰ!E[�z��m�Nq���-vQ%'N&na�F5��>h{�, vm{��ގu=��� o���-��v@�i|�iߖ�=�v�O�|0�y�v�x\�C���^-G�����8�˰������!%�z1kF�4;��ʯ�-�=��qؗ���K�)]��
M;U��Ѷ�Z�E���L>�o�7`���3!��|%[sZ�~�Yh!f�A�� Ǝ+m�M�����篾Y��qĈo�i��e�&@�Q�i)�O^��G&i:M �.ϔIN��YWz�$���U��i���#:T3۰]o�e}��������-{���2���1*�r������D��Q�����Ʒ��r q>�Ƙ���d�o��ܐT�Ӳ:5$,#�����Ƞbi'%H��;cT�G�N����HW�J�9Ye��X�[��DN���*�9�*s��^���A�d�-	\� ��7���2�X���;�pq[,���I6~�e�	Gc}����fМ�3���^����:�e/�$*�:�]��d�J�P���W����&�8!��'4�A��2T�pf������E�R@�K,��.�q�6�)Qq��ڝ�NJ��5���j�h-{���%���3R��G��}$�g��~��a��yC:�s�rB&�B	�YV�mz��� �����I�^�s���y�z�LR��$���D!��LW;���Tz&�3_�w�!��0�I��R�×1|�PNA��!K��P�ILg�WM�Pa\솖�oj|����j�����qjI�J6|6g�T���F��{(q��g8A�ݐUQ}t>B����`��W2��J��j��k��E3�0�o1�ӽ�;2@��]����ԣ_J�9v���R������اݿ�R�Khs�N0���p��jo����h,*�����Am9T,,�f3�P�ʿ\	-�jc� C�i����*�bg���z�-:�O��0�Wb
�W�Ӯ���)��p�4b����y��`�����ͥ�J�׶�$t��(5(:�6j��%Wz|w&�4�z��C�� �~��Lv�03��e���H�b����Ϡ�܆�:>
�N�3P��#䨐7)�J�Ӫ�\�zȌ��d����n�E��`9�����.$��~-PڦY������K�J��@L���o�����L�V�̃��41����r(�o*v�eL��8T�'�s=���:A��Y���b,���̋Ha��S���B��}b�><&Q�&ƨ�v���]���pEac_40�Lf꒶z!/���œޛm���6֏ � V�)�%�}�8�6<4��k0	*\����ڰ4`"Ͼ\,)C��^�*�'K�]���j�]&�ǈ2�e�-�<� �}J�o)��X��*�?j̙�T�k��R����}uj-�z����U��7~4�;qթ�4L�1$p<