XlxV64EB    5cc8    1430�ݥ��.�Rʅ�T^���S��͡Q�h"��r�ȫ��H(�MH�c%��~jPg�W��/� ���v�<���Q���{Z,6�1f6,Ʈ�����RH�"�\�f��B�j����ݡ0~l����� y����q�4����'� v�4���t��]aJ�vP���[6@_�A6��HX���<5�(�eY����c��d�9Mg[��@�d����K�"�iK��dj��(������jȠ�]�H�.]��<�#�bc�-B�=�h	p��>�� �9�f��� #����?��z��]h^w\:f�����G0PE}���P����C�'�kq�Қ��.6�K��
���>�ChmL>���c�]�ސ���a����ԯl�I�U�<�O��~��Ò��EE�p�����׭�&��HIL��`T���9x,��Q��&e�6���e���X�5�W���m�����[���R�z�o�������W���M����3&� �F����e]�Ӫ՛�?����g��KԒֲ��dUYY�A�$Xи̏�	P�)��߃�[�Ƞ?�,Q�|��-���tDd�Z`P�Uk���h�,�:��ôy�P��@?����d@�LI�K��K(3����s0V!>e��!�5TE��
!Q1X��	�>��gș} ��@NU���L���7��{�p�f���r��#8G�%�:�+��L΢aG.u�c�H�� 4����3N�Cd���;D~��a�)h�����W>d�ri�$l���O�hΊM�բ�F����[ ��T�l�ߙ�X.Yc1u�+�~�e%tSҟ�D
�[�F0Jq����%ϵn3;[O��:��o�Hډ�-���������qZ��G7��ƀ��'^׵�2�^�[��.rk%#a0xC��=�r�y���<th�+��&7�@DM��Z��1�`R��p��UQ>P짳Է����Ք` U���<����<r�!�����a���)^�o}9`=R7���_%7�=+�{��n ysŎ��W�F��3�k���B^|�[�o?������I��t»+�ܴ���<�m�2'���t�����M�7z�QV
�i�%l�@ǒ�6u2$�D������Ƙ*}u^T�͠��<���ȧ��h��NU��dt�L���7<�aಹXu�7'+I>�y�y��!a@iQ?x\,o�	%!����A���Zr������Ѕ�I���Rѭ��?�R=@e��w}n�:����VM쭧@�:N(o.`�屲_��<Â����u�X�_y6�yWׯ�y�Lz"�9�l8I��#�Dp61��5������V�!��Z΀܂ ��Ii�MFۺ�+��5��i�Yk�V��Pl
2�y��v�[�(�>���5M�M3n¼
5GVcs���:U<��uݱ��S1����D��"��\��Ty�KE�)����bƦ*v��`4�(�(���%�Q�E��-��N�`9W�	ِe��^�y��n��B�;�JC�R5���TO���x�Q��OvN$d��j���tT�^?K�_��u�����m�]Ga/6Lg���诂4�w��Pj�q���rR�	ԹEJ�8$Y\����8�[&���QS�mc��칁��8�$�t�,dh9�/#�v]_�.��4�H�H�?KT�ڏ�B3��F�Oi?;�,ȐM���j�Rh��ˆmJ���^�<�~��먛���8V����}�����[�%_z���?�Ӎv0$";��O|-����9��lڅ=�b�k�I����p�I��a����h��ُ�!0<Z���8�#��̵mwV�B��� ��g�䆩�Wg Z�LCR[4*Z�O.m��ZuKK��k�aR�Ul5��g�'d-��0Y���_�~- Ⓞ����<W�$�f2��L�y� d	�@a��ln�ۈ7��K�b���������F����(v���%��o�9IZg"{�>���Ɠ/d���f��M�U+j%JO��v�ᵠ;aHII�wџ��p��7��
H��O�^���ATθ�ɥ��"޹˼p+���*����D�����V�}���0/T�J��W�����DvZ�0�+�����PѰi�z����+6C��<��Z�3΋�{�Á�>��!�ь�O|f�:2�P<��SlL�Ta@��F
��
f
H�*� �5�����!
�Wq�
O�|�wD�#91��Le2	ze�o���R��\�QS^�׌���5ө:��Fwք_:�4)�f5-�=;Oנ�MQ�bU 
x˓��s=�����l!	��9!��C����h&b
�J���c�H�e���{�D�d��E��q���O�����B�h��J#��G��8i�Ӡ	�f�9Ӻ� (a���I������<��Ep��Xm�j.��s�����C^�K���[H院W�F��p9V;�E�Dpc�N����ӮW����!V�0�\#�(ֶ���nBZ�梙�]»b^���U�[�=����yB7\sv��;{%�����n#M�\O�u�nNh���K�	��7.+�h�	%�!�Ħ�b�aR6q�H/<�R�}�<Ps:���Ԉ�� x�[� �%ʲ�$hm�����R�~��Qe�ѺVuJѺI��L�$F0����ȩ$ ��fj:���0P�=9�=�Ƀ�Ŭ�Lt�a"�8k �M��wzmX����\4���ieʫ��Љ��W�D���c�E �I��� ,n�7���s�5�y@���w��a�˱��Mv��%n�Ϋ�'�O�jP�+��ivs��]�S��{�9�AF��/a�����kR���f|�O���.���E0�7	�y��d����~RUe�]�p�T::��w�t�V��+F�!�q}cr�Wt��� �4������C�;�;&�d�ȡ�����f��k�J�@qw0bM�J�6�?l��OM�s�v�>+�U��yF�D/��w�\�c �����(�5���j>����ڤo�C�w�ؐc����m��J����ɪ�џ�p���v�P��z��rs�7�`��Y�LU
}Bھ;���B�Px0;�ـSfW�[��`�O�A��Oj�+�"Ζ�P�7 �5�|M+��/�׮��y@�^�[g�M?��&����䂂|��[̀[*�ײVF׵M�q�\۵T.MC輏+g
�Ј0�&����4Z��i����\|bY�<AT>��ehLE�lI7�>��l���z��>�c�<��i��t��cz�X�H�B�flÑ�rC�Nw���T B��џXxS����?�-�qG)@�J��%�Mh��,,�"p
A�E,
��� :X봈�.6۲K��O�_r�.����!���l�N+t��سǅ��؉�64�l!�<�x��ܕ۴P���1uE9��5KG4
)d�t��k�
�d�o�8���j�F���q������T��Cq�q=��fImpK��tu��y��)�L��qf��=�C|�C�m|!�P%u��"���]9o��ԫj� ������@?��8����"��~v{'��*�j`�r. �u:!���N�8q��x��Dmqe��.2��
7��r|Ft]}��v�P�P(�,�ݖ,˭��au���<�,+��ȿCKr��QK�N�o�m��;�O���G:��'��mh�^߿�~	��E&G�^��<�� ���n쥿�U&s̊Hr���-ڙJG
T��c����dȟ[�V���0���/��YY/&�zߨ�rE��@%�jޮ�6|�fd �h�<VN�$l�7XQ���W���+$ӓ�۝_(Iջ.D��-�ƪ���7ݶ	�&��ٜl����a�h������	�ϛ�#�ڣO9t�a���O�e�Ef�.6�-��[}����*ku02�Cx4�$F��IBܙ&��cq��Ԃ��~���A05�?���Yٿ�߇�J/u��n�ξHn0�թ��+l���@�\�\~j�^�(��CyE_��HP [�<v��7/����O����k�ߺ�,�;]��/c���L��x^�6#��v�Ṓ�:i�q�O��A����#���y@wX�n�sR�È��V�[��Z�"L���/05���W��e/x_���F��/���$�\���V%Bn�D}޸	�dڰ�}/�ņG�[fλG���&I����@��f�=�;`�g�o��:�f4Z��/�8t�a����8�ŧ��Q��B��[�B�P��ux���H64��GY�?��܊��Wr(+n+��J�d&��箸����0aڭDq6�F�<�q��Vr�bÍk��)`����5cx����jΗ����T�zЀ��>&O[�@V���\��fa�r����ħ�'�-�5-�+�]"DiWq���r�X���Kݿ����p#F`��.��V�����9}�紏���.�<(����e:f�C|����+�����Z����ƀ4�t��K�n@�rc'�4���>/�7X!�b���&�Y���O"ݦA<��˜�w&h�y�%��#�o�2q�.	�@��Д��W�G�̨(���?��W��1�Au��E\V����c>D�k��.]��׾,��ldqM���������MɑE�ὲEN~Y8�L˴p
{iB3�4s��6@
��5rZ�������t�So_�t��G�8�an�A)� �/�F�*��(���G����\�,����m��o�e!x��U��g�/���.�B�>O~h��G�^� .�v�G�pw���D���)��"!���K���L�Y��Iboy��:�yQ��̻A~O}T�
�����J�uokPV�A���{�O���L�����8/tZ��?�6_/�):51/�p}e�� �:���:	��:��H�T'�i����(5`\y��(ڍ$&f�^��2e0����T��n��F���甑�r2$� lJ�z$M�}qT%�5�8�!��<�z�χ q� _���#w|r�����V�����c�c��b�[2	� ��;��tc�덺|#R���_�."�	���E��d1�b���ҷ�u�ܣrX�5љ?��(b��{DT���s6�,]�Лj�S���e�E��