XlxV64EB    2e17     d30�[�7��D �ߚk�y���^�Ŕ�ܦ�_,{�g��*�t��G��U���E��cvoC�����d�]◺�މi��c���bJ{�ac�ʎ��N������A�ɰ��i5�00�5�4��$S=�Ӥ������=!���WXYc�Ō�Y�+��Vp��p��"���Ә#�5g8R�e,�� 1S�k��e��l�Il�b�=��0��;T	YЪ���ݝ�w�s�<�pu(�\n伦��?�M��$w�b���:f��k�$�+}���D\34(	���І#�g̵��π�����z��|��C��[��
���9� �`[�>Ķv���IdR��(���ȡ1�_�)8X)�&�Ae.�{��N�U~+lz(����.ȗ�*x���[��xN�ɝ��k�6�/oq1��_������A[�I�#��-"R#L��Y���,Y�b��qOdǜ&�!��	��ķ�V���ǹ��x�o�F�Ⴠ�xz}��J@/�(;Uu@�y5^��u���tX�$�+X=nEś���K�ѱ�F�HB��<@����Fz-���)�|BV�E�F�Fan �^!�ڟ��R��?�C��]��L�})V L4�V7�����d/�Nj`߻�>��/��7��g�Q%��x0���Xۚ�W��4M�#����R.�
�LR�Mm�e����יW�v*�!��.�2u�,s��[�(�Ӭ�}��IN;��	G%^�����h�zN��Z�*\w�k�>ަ�[���T�sv����L�Ŧ����!�P���.\)/���Lf4�T�[o���l���.���"T�~F6�w������n������M�i��=a�Bi�~��a۲�ú<���p�;͠��x0(���C!�Z7���S
�3XH����0�|��y�*؆��k������W9yc���#�8�r�����
~d����x+�2l��Ԭ�������%�#�n���b������5g���y��]�6��^��4�T�%�� �v��V����P�7�u�+�9�u��a��Up6ov"��TZV�������$��>o�ήY��i��^�8�$G{��<�	 gj�޶��E���罥�ꗚ����iZ2_��U~��}uxUy	<��je��Q�M��(q���E$��8�\5���ۥ�����q��jľ�ymhfN��1�Y>�y�v�"�p�濼 ԥ��)I��[��P��e�O���I����Z�JoS���8ㄅ}V&���IKad
>�#�
��z[�ɬ���\gj�l��P�����3Q9	�{��k$�a��*�1n����7�&_Q�Ӹ�p�`�y��y�\Fݎ����]�y����]F>s�e{h�'���(�E������kJtY|��i��%EAHz@#�:��t1���)W�nYM��#+(<K��S��B۶�d-,�|�m0�ʋq�~�d�B�,�;F�T��tBNΗ�%M�u�8�f��D���k:�� {�f���� �c"�S�e�}�*>����0���$��޵�
l��0�"^zW�.6\�H�m�*W����P����9W��+�
N�>�C�$��̃�"#�f�3y��	��%n�����UHJO��G�Q��O"'��c�G5Kx�ٲ��h�HhQ�l�	U���=s_�Uƌ����M�Z� ���V��^_�º���V��e����
Y�)F�Y�nW����/.+'7���[|S/.{�F���Ւ���L���k�l��m�@D2);�r9il��J���d�D�?%��'�<�|V4�:͔?M�uX<Y�}�,�d#�� ��f�-���V�QS1�e~����lW�]�W'�鼿���6D��Ob�C�KK7p`S�Ƕz�Dq������/�{�pnQD���!�����@v���3,��>��(�H���ӎ~�p�DȎ(�Cv ��O��u�yT�����8�Wn�n����Qڠ���qZ���xy)3�� �y��ź�ya@��J�����T� т�;���rA�`��~A_��H}�sf�.*�$w�b�=����2��Br��	�F�̚T}�Y!8��=�髗��YR/�؅��4�1V�#CQ<�0�p�5~�V�F�8�H��a�ͪV����x;>#Nn9B��#�,.ge8��v�&+�<}T�EnEH���2��0 J-M�R�-OVj魳@�c2�9�_��?��9�}�094!S??o���5�h�LOp
�
%�X�p�C��y��x�V<8qȩ�_�p� �����c�����&��;�zILA������'q%�c�|�e}t�X�Z1'ts}xy �``�G��?��+�{��
���"���BI�*T�׋����z?4�0�wq�q���q�|��,�PI�e��æ��0��߅m{�l��'�/4g�7K䣸�n�'Y!��,P�\��p QƆ�/�2,ʘ�9�#�g�r��t<=��]���$��b���z�<��_d��I4��8�;��:5�m�V���&��øŢ��#S�1��D�)��4>���G�7�_�~P  xu}Ek>��C�ktmu���ދ���'���w�i���l9��Y̸Br9��F|9R�������|����r�Ѧ]n8�-��Q7�\�)َ��R��F�/X���� h݉��˽�m1����#���9��T2��J����n�l@�?����}Я�k�<ȏ։҉>Q�̦$�n�ӎ�	�G���.������>S��bN��5��n0V�=�*��i&�Qi���p��
���Tӝ@��W#�߹zp7#%7�;�8f�����\p��8�,_B3������n�V��u��7,;��8Q���� <��T��h;�2-�Dg�I���csQ{���<6�P�^A�p�{����3g������kIw_ �F�h��R����M�ɣ!_O����.���<�_�*,#�bƪ�T Θ�H�MF|;y��j�eSti;�Y��Hӷ�;� �eF5&�M1���_�����
��y����ֻB1y�3�b�����Y�����싀����!�`���R�*Tm�� ��_�dr
[>d���.����bb�/j-*�������h���<�E���X�nϔQ'6� }��9_!'_ɁӒ|-˙�œUfr9��Q���ԑ�!�9�%���A��-�:@mZ[nyq��x��cȆ~[MםW�-�W�p�l�����H���"C�.�qKw���p���B@��2]2 e)ƕ�Y�LO6����s�^��\l�f���;���'x�T�Q���e���0�oy�e�\6�� W}�P]d�lAl�����(\