XlxV64EB    73ed    1710�+9���!g��r�M��ړ����i�#8��{���
��}8{)�[a��)���M�8�J��WY:�I =w�>��k+6#�q�PK}�\��f|5�]}=7[N�Σ4�A�L�LD��(X��������*���ȷ�a��XpH$�(]���C�aqo�m��g a��ɝ��E���L�g6��yD
��ʁ1����U��1'q�J�*�Mp��!��J��ƿ&�_2�b�jH+�w^��ደ{g::&n����g)��WŻ6��]E�Ս;����ӎs��-���G:�Q�>�HL�.X�0���r��.7�	T����ďˏ)�	���u3�[�O}�G��q����n��P����ܬ�08n�j=�ŧL���&&�w�FI Be�q˚G���˕�접�1�d���e(����#)�$ױ=_̦3�f2`������(r�3���	��$n!���8���ܧ��#F	�F�$�����-W
Lv�x� �=���R�Vh��p��[ם��k�g��Ǘ�7��+��dI�
g��_�Y�
��'�a�2T��>��[�ޕ���a����}�[*������x�U��x�';v�ve��`3i���4�8g&uw޳�qCީ��޸�c����h�4%������5��q1A�d�BM�_lj(4�e�!6mt�;*�M���ek���1~#uz��cm{+�4ͨ�̭J��YO�|�'�H!5$�E�]e�k�q%_Zש�`�G j�}���;\�-]�B����$�X���De���f0ʑ�EF�6���pqpߊf�0��	���A���������7O¡�	F#�`3^��qqLL@�;�F�6���$l���+�3�	,]�k��q�hL��Rn!>ֻw$V�j�Tt�ӏ��g\N%x0	y:"� �*I7X�����x1�#>�N�Ni�7'�4�\��l 	��_;q���쉷���Ԫ�sѡ��������P�f�ݨ�TlA5p��HW�s�������گ�I4�Z��C[�oY��!`�y�rՎ�?�VP�E�ad�!<3�:���L+� +n�p~ 1�%�<�τ�'"B�A��^�"����>}8x:�P�?��ZH�^��Na��h
y}�n:�B���Z>��@��O����+���4��r^����
v2� ���ػ�l�ņ�j�1�1�L�T�:=3��p,�>Z���P����4�u���I/Y�_5�<��%9Oh�;�nl߁7��)��C�{�J��/�H
������74�RQn����ƴ������b �nh��+��,p�cL[y�tٖ�/hK��C�&�-X�J�?�,�"pyL�!�՟���Z�=l��K�xyڼH��U	7N�������5ȭ��C"�t��Tв3/�>��~��c�Bu[}Q��I ���H�o��Y���i���;l]��H�E��7t��p'z���p��P�d�1j�T�n�jR��S�_z��wC`YP��NQ"\&�?t�����i��X#j�3�:G�)�Al���ÐE��$k��gEJ�x8������~O��GV�X��׽�`���oqҮ�#���BSЯ���Ix���C�T���³aTh�0������λ����j�3M�k�����i�&o��m�}�%⏦#�~$��I���wڷ�o��eE~�:��S�q@o��ĥt��i{�?���s�W?o]�B��q�#��fT���F����:�#��&T�~��p3�+�K��8�Y�D3sr:��n�&'�G�M��4��-�J��C D�R�M[_V��V�\L���T��7��Б�kd�s���	=�Z�j���omo�?���-�qG��M�C��n��A$�7��w�ђ��W�pؿ7��d.~v�ϸ��^�T��3�8�ޅ<�fXZ�i�`������+�M��~C���k�����S�&`��H'T�j�V�<�vg�!RO*�h�R�$T����D����L���Pg?s�\�G�0S��e@L���w4���ʝ���VŮʽ
��<m`�n� &���Ƌ�M�W�5�! �z���Wo\ �樂�X���E�1�E춲�R�h�~J1����B��)��x��숌e�O�̓��Ò��/<�\��ߒa�b��i}3���yo{��?kG����6OQ��5�Y�lzY�RU]Z���'5m��m������o�&]�F͂��Y�!�.>�7ѫ�Y%NF@~����1 ��L]pQ%U��U4:�����(u�!jZ-h�(�4I���_��v���z��z]r|�.�Vq�dh�������I��kY��^���Zj?}��ԥ�R�Rl�z��f���M�X7���C`�$uK���)���H��3�{�Df<;gU�Z�I�|� ,�V?hR�i)f�z�zፊ�AW-�I8,��^��u �Zr�����H)���V����j�q>�I@����s?�y����\E��XeI	%
�ׇ��z�7?}��1hQ9G�2H5�nയ���>��;8��<1�b*9-���j2�LIUe'������y��@g������a���o7�8(,X��-��wZON���h�t���(�����!)���Q�]��;~����#f�{�F��g��D��w��c{W1���3�@�Tf�~�/#(�uYbKY�F�Z�{?���<��=v[i3��>U��dL���t�My:����ފg��dQ"y�̺������-�vĐb�R�@5��{J4�0d�'e�Sc�)���*&�{ĸ|/cA��R��_�ZR��.w�!��ׇZ�FXS�!"e~/�ɩA ��;R7I���x��6�u�`�fN�Gf�"Qrd�8�.�(-PiWoA!R�Us�ĝ!^ruC�*mS��O;F�f�_�h��Ft��H��slRu�P��t%�a���9,�6�p��9�T��9�me���p�}^~�����J1�4���k��D���
!���/�F\�{RƉ������U��s�9�|`��=�ꎧF-w;�F�.�cJp���뢮*�5�E2k���n=]�C���[��0��fOJ�_�
Zo�"�W|jx�q�G<{j���:F՘�yh�k��-Y�0�l�ȷ�d'L�Y���6z��&F����V#���Za��	�&vTG":s�]o�}�Aa�3*ΒP�m�@����q��?;�f�&H��8;�FgR@�03e7��?>��)3��5�A(��qR��!���W�;U�|� �6H�a�#��*k
�f^� `�j��v�� ��}�#e'������㳣�����LdD�m	R$J�{�hG,)Aaz�'�h�K��U��D=/�AlӽU�B��]���3�H4��ޘε(m�������C7.Y���,�bm�Tk��k�n~r�X�^TZ3����'g��#c�-�	,�`���U���yq/L�9"�=�=�<�w3G�T�h??�`΂w�S�+��БG�T��K"�/����i, J�9RZ��`o�N-�3���|[�c,�j*�ڿ�!��*�+kT�}j�\�.�7��ʞ@3nĢA���$�ĦY &s�V�j�?�Rn0 �ѩ�|�̊؍M:^:�-SF����7m� �	��©i�ښ�yh���&D�XP?�;N��l��>M��ϛé6Y`�N����ۤV�ɘ-K�=T��W��T�m�ֈU�g���z�rexL�p뾴�I�z�[�[�12(���5Ԧ��+MQ?]+W~亮`��-Tc\%�j���2������?3�7����ş�5�뙈yoH�y�����Y��K�x�NOJ�}�@���5gV��$\������v�rlʮ�f1gW�ڂ�f�'�q@?>��P���--w�R�d�`E�:�ؤ���	R�=������tr2yoGi��z�����V��	���/Ue����]=���q*��=��P���HيROR�CfpR��ì��D䦼��SZ���S������J^��Ha���{oq��;"f>�ֻR��4��?�J�	%���{z��^i���i?�vN�YR*��"�%c~�I���ȋ�qU�ƞ����-V��X�N�,�:�M,���(�r2I�%���<�¥VV��?7IY���AչG��;�����#����E�T\�U?�������_���*hLn�X���4Y"*Y.2�i$bk��)�ŚA��DA�yWe�n��**��m�S���u��-��8M!2�S"y��d���״p60���=�ѣ�2�H��焔�/�g�x����lvW�	���[��~�mDG,`�ds��1�"��:!SY3���~E��+Qk$���ݱr�Fn��TI�4]��m�F��#�8����VMK� �믯�%\�'��	���9�͡�
��F.���Y�O��m�O�C����z�j�S�2x�y1���*	$R7\~ĸ_���|������Mv��`���A�T|�S��h��;S�@	 h�]M�6`�5�5.<��ꮴ�_�?|!	�*
���J�j����G̤֜���p����,ױ��{�nv�h������Ĝץ�M�ݞ*-�wJ��2��(`\������yePQօlK|[Hr�|�j�F�TqcM��[����`���t���Lt����}��#����:5|�9'qOʮ��d��+x�"7���O*OO�Ҿ��'�2��N�����ݸ���w:��	|d�ط� ���޾!n���	M�Ir���jwk���娴A�|h��T+U�I=+���ض��D�.�������U}LA2��	�)+�龿�1v�4i`���}M!�:�.	�Jp ts�y|mN�䪥�(<�V�ƍC�ע�l�����{�.��C����#ʣ��KB5\<�&H���bn��'6/>x˶]�F��/-��+ %����|+�\�b��I�Q���D����KUT�%��G�;��]�d}��&�.�0�L�xv��{Z �H�|�M������x�{*H��t��+Ďko�T��2����#q���N�G�k �{�,���;��7ʾ`�����GjaT�T�3a���1�P��y�e����r��}�;��������Qv-X�A�7͟�D�i�1��Q �?��+*-�:��(G�"Ǖ~V���]���T�U���Q�Vzd��y�>"����XJL�]/ń��J��D��#Z{���^�	�2�ta���ؙ ���~(�;�����.��'=���td!��/�/�?o���"�dGⓨ�SExm�50z�N2�v-~\���/@ل�U�''l%�"��,R�,s�#�\U�,
!���1�O�%�`+d%>���՝J|B�]�I�Ss��@��R���,&,=���~����8�-�X.)��
�rd�	�)�@��/xPڇ����M��P� ��<�3d���J�8+�'U�dǼH�8�o��^�������xJ�q��m�>:c�@/P��E�;zn7��b��p\#,�fT�V-�M����
��N�<��B����
�"ǂJ�A�	��8�=�Ȯ�HƂU�W��ö��������cZiKK�]�ǚܡ7��?g����о�0����qd�q���G���T;�o�BQ5W����������|Hm�;�=��� ��) n������e��g9�A9��"�L�"}Q��댷���$Z�y>H�����.��*t����/jX��V������R�g��*�a�~'����~�Dz{4V�}�?e9���S�&'$ɹ1DUO�;��-QW���n}W���kU�'6Ut�i�dEcw��ӳ�>�