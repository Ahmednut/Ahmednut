XlxV64EB    191e     9b0����n
ղ�Z���a�t�/�XN��~mcV�~��5����RƄ�ȵ����K�W/��W�6�Pîn��\��q�.�n���!z�_	�`���k�U���*��B���t��z�_иfŁ~�|@VЂ�O1�j�0���ɿת˥�e�DҖr|b���OW�R)�+n���Az��1�"�JP5�@"�;Q}�{�����٨ٰ��6�Sӗ��3����{�SJ���3} ���������>t\��� � �a�D9���˰��#�`jR	��k�?�.�R=�ܩ��3��fˬ�dŇ�Z��(,5�i/j|��#CW|��$����Q,�Y7O�X�s�uジ��?��y`[Ў1�x��#�ڥ�K1ڨ������.�	�m�,�C��R�����r>)������twu���M&(�+����s�O��.x�8��3�h���^��#����>�׬Y��OH��Vu`U�r��c� ��SZHD���͔Ϗ��=��P�-��������;Y������6Q'���1�-k��
J7�-��E�*]����;i�YҔ�k�Ud�����Ik���ꣻ�=�m8���<-G�`�ml��0��-r�D<�K��7���ڐD:�Mg��v����k=��=xh�ROB��� ����/��dr�>��sb�w>G�	���C�3Y������%�E�?^6K{xF.Cq�9�vr�L��� ��7nXi��wȺ���m7��7,�3LX����V�\�)c�7v9�k�ئ[��0V�4 ���V�M8-g����9��1�5�;�,�\��"�&���o���6�xE�sX��X���.p��H?q P�UA��hh�g�e��Y��A��TU�0ɿ������WTw7n�w���_�RpH��3��ID�W���D��Ͼ�h�2�$�Gn�����M�A�q�D�zS���D��_|�w�6���<Z#Os�MuŢ�G��9����D�D����}���*S�֝�N���?���b�Bg���|�6������/)6w���CE	��z�~�{ܱ_N��@��H�5��fh7�s)�"CMp�aw)"Źl`�N�ݍu�*q!<ʤmR����ؼw_Ly����(�+pEo@�mS����ڴМܽ(��1�򥪸���m�i8�܎A�Ep���e[�Z�b �C���}��`����5�lB!�락��r��Y�|�?|S�]�e��������9��̗!(Y����đOJr��}�js��ud�|J���`>�Xc}t���rx�Ё�c��{{�Yn�R&F��?�k� �	��Bм�%dx�v{�$��{*�CLdB�Ԟ!���`A\S��vrF����r�$��i�&P��k�c]�(�����v�L彲O ��vWt���9���ݻY����̸0�s��[���@�F%"�t��
AY�1Y]l���.]�����|�top9O���>y�e"�C
�#鄅~�@F�$g�
*n���T��ڂ>\!�C��ph|m�]�I$���w�p�X���6�,���	�V&@)�,jWr>��#",E�D��`���cy|��EBGY(�P*rs�d�Ĳ�v	伅>ke@f��?�g���7�z�L��Uˊ�2<��@���B���:d��
8CX8!�
>��pX��>�D-�Ź�g���mrQ�a�H�M�^�Xw�Y�U�Q�E���<��8�3ҐFF�w(�=�>=O���%,)ԸC<��c�0�~K�$QL��c�k��-��z�yޘ�^r�@�F�NdjEP?4�a��H��%�;���1�X@N�}����t����<i25��ODޏ�@w	��:�)��Y�� Zh��3v��3��^9N��խ��u$�.ڐ�C��XS�N>S��G���Q-f��K��54al�B�.���@ؠ�?��)k�!̅4�z�є�i��C��f�w��9�����d!��6}a��L�C�!���y�)�A�%]!λn���M�/u��/`4���z �C�8��DO�,��v��k�Ȏ٢{v6<���&x��r��cv�QLD9Z��mI���x��߂�T��Ȋ<���C��6���0n�]��c���S}�� ��O
C��ż�h.�1sYy�s'
-�!�Խ���fϓdq��֤��s�j��
<R+��6����p�B2�H�yY�},�5��ov�|�������ށr�.ɷZ��y/O�TH?gw #�¿	�/�G�%Q������YX��� 2k�m�t�g���e�Ź��4���ٲ���'�F�� {m��e�ǩRk�`E��".�|�I4m����B)������( �4�"��8�#9L�%2��ӔL��(_��m*���iv�-�n��WȮ��8�m1�{�)Z;�x�P� f�
����£7|4*nʢ%�Q~��hj%lmQ�3�;t�5�ٟ�/(o���*�:I