XlxV64EB    fa00    2f70稁	db���=�5�	q Pk�`Vɨ8��P���+��!g���J	
&��Y|l"p9�O�~C�իg o����2]����'�Y��>�k�������@����A�|����Q �&x9?�fB� n���n}��mb��l��hPkQ,�o��A0�oy��;}0�9�����-�[��t�į�A^�t���'�g�<��5��.Nĩ��՗����s��+�:�Rry���j^[��>�lqڥ���z��W�4�;���W�s�$�M��]��[��Q�O���P��L>�V�G���۲��'+���8$g�X�j<���:NtMH �,��x|�!�D���=�.9��Ǖ ��X����N}=�}Ny��wga)�7*-z�U9�e��mL�����a��e���0�w�
�l,��*Tǲ�F+O]h�px�+��v��̗�sn�<�Q�I�|���0�O�V���l6��L����%_H�4h"��J�g�E��!Qu'��f����N,�<?��˘v35{�Z�0m����3���=n$hJ�����ܩ�A��"�d���5����3>�hZ�.Y;!�ۚT9	hm����.����K�3c�S�gEI�/MA=��" ��\s�7��c����F�c�X�Z.u�ar�XI�o�����ß�}�9��O&x���j�su�\���
��ɇK�!Z�$x��$t�Ev{xW~4ж��1m�[�P��Z��[�@���7ʁ"D$1��r���Ӂ��Yd�G������:���~�9���Ò��J����Ė%��%T��ε�~T$�72�}'F�SSIR����Y7�>�k-����=*}����+��p�fiJ���D k�e�������<{tHO����Qq�q��9�L6�m�~C�ʇ��>��Iy��{	�n�Lbl��.�d�>���E��2�%�؝ue=P)q���c�s���$_J�I�]�%��	�+#�o)O���ˍd�p�S���d�>�97H�L����A�4I$����>y�%eH�!�J���!z���)�*�#mDg��jy���O�f���Ke�I��a����(�o�����}�Q�9kP; A��W���5kZ
��ah3�{�i�=�p�3S�!h�*s]�|�P$���ѵ��Bi����I)�-['(��sՠ���+�l���E{e�.�sؽ��76�uLa4���m��+�^���Ga���)�/�Le7�>ܒ)��b���e�Lsu��ީ��ع�M=��*VO�+�:ohz�� u�O�`o��
|*@�Z�Ps����i�|�u�?��?�H�+}u�gW�Ӂ������m��a1T=��k?��q���M�;�<����b�y�E�C�<�>�<Guo�1q���o�!�W*�s�%��Q�l�#�����ӕIU��KǕ���d��"׭
(5�yЗ�m"���ݯړ8����IG�MO���>ƅM^��M;�`0���.cW�+�/����S�p�&rvRXF�Ej��J!�ς�.Hz7?p�Ԙ=�=@�}�	�|�^^����n�Y����$D���T��0h�����d�����6��A�P�V��Eާ�,��ՔX(@��b��ƾ�t��"��l���L�AY����Q�~��ޮ�w�e^�-���6�8 ʗC䤍�N���&�ު����s���CVS�Z�Q4�@��X�TK%�-L�6��<
��t�X�b��s��R���:NOm�N<�N�}'i<�����b;R�>S�7�h��W�E��!�g9YU�X͜k���W���[`��Xc
���7c��E�w�.l�D,fo;�\����bH+p=xjld��ם���Ӂ�
);���u�9 $5�I5M!�>@3������(b��o�T�Od�		_�R�����@|���SͲb���%n�G�[3ZCw���/x�Eg�x������l�@\w?1�q)�u�\�>*u{��<;�@����շ��M�̫�:�A���Ϸ�aA\�9_8������a��*��ng����"�z�I��	-�I/L�k�/s�ۖt������*a���ժ�o 1
�^4��ֽN��:���3/�(֋E�X�W�}!*���	�u&]�o�c�
� lF^�/b�r,;���� ������pƤ��k��q���Ȁr�#�5��Q�əB�3{� ��`�ӱl4��� =�I�g.��nN�!�R�֐��a*#ĉ���Guq�Vcډ��boI�l(r�m ��%��LA�!�l��N;��=e���3�D?�ZH�l�m�0��=m�`��rU0�:? �7|�pH��	\�y}ꆬ�hV�%v0�X+���=�������c�n����������9a�İ�М�]=._,���X�n�q��v�}Uw�^n-��H<X�2R�$�B�Ğ�g�$J<�D�ǭ�Rk�A+5��;]!hJ�����190�mR�ٺ�)qd�?`��PZ�u�۫���fМ�^(��n.[z�:Ŏ!E�	��?\@�b�I
X��&�RX�̮J��a���6�
zs}��=��ƤF�υ�����/OКO�"�Wq�3���z����Bb�=�y�dRgJR��ԩ^�A��4�����6���3�ʠ�a�IF��qoPϹF�%E��/�~��uzK5O��:�n��mX�H�8�bK�ܵP9��t���92N�v-��18���E/����	,s#��|��b�){�T{����L�)��CL�rC�N��lX
�v������ٟ�
=�<�nb��UG�R�ضC�&�3���&�bc��N�l��/�rYw`!�t�������dF���F��X�',�r;ޜ�&8[Vr)j�'�A|O*Q�󣶬�79
b�Dia7�x��Q�-;�g���~�e����n0?ՕmmONV�<��Q��z���)���<���oi{�{�{c�͍������.t�I�B{h��W\G��l�@8u�u��wM��fx��j���gτ��})T o�OW���Ri�������Eis@ްͺ�.�k���s��dp+9kH�ޭ�ey܋�v�%=ȭ�t�S-��~U�'p�x��iS}��%����i���~�ef_�CD�jdD�ܶ�^!�y v<�!^�|C*G�$4�GE�9�c�W4Lk��^!:�˕��Щ?mmm�P�y���Hл�4#L��3���A{Dk�AY��V�����7����B�3�GX�ګ���E"dF��a�	D���[��yo� i������'�MΖ���3�)w�G�3F ��_~Z�m>eJ����^}x����TXP"�&(d�)��L*EtWd����E)���uH>��Pd��1D���K�s�Y[6�� �.Tߗ�������
�*Y���I�w���&Ԭ%�����Uj���h,��2�z�B�o�L�t$���2/ȩ��0�v�d�� LA�QY揋k}xOV�y�@g\�=;u�ŵ�R�cǗf�lPl��Nn;� g⸪�
cö�WT}�f ��-Ʒ�?L��():������4Q�"��	o��O�6��75GDF�[���L�݌��Գ��fu�b��zX&�L��J�N�L1��H�]�0�v�s�n��	���? g>k j%�Z����_�Q�е�;�������
\U.�\Ϭc�q�Q��#cc���iG���pb�� ��"S�`z�hu�s�Q�H��<Rn~m3�+����?oB�������Q��,�E���c�������i!t M�@��r���G�Rh���T�RDq�sk�P��t
ve'�'����)��/�w+r�g�D��������x��;U���5=A�t;��K&��pv�=�t�i�+ �
�6Ó`vh�pK�z�m��5���J���~���W�$B,���p���D���߽� ���������(%˩�B!�V$~٦9 iԎ�� �4��P��6˞,%����D�ù��f�w�7h7���>w�N`��ϳ�&�V,��g��ĵv?�S��� +.AO��r�!70T�?&��(ޒǎV;�]�V��e%p�����4�Ǜ���@�p��N�ax�g�Gh;�ܟLC[�� xhZ�t��C�)<w� DK�a!%��y�X+s}?�b��cJ�k	�J�a"�[����\B�����n�H����< ����j*r���q��������BHC}��s�sT�z�cR`J+��V�m�s���#�49�7
OU�/a���J*�U<.�^&���������%'��K:��<�|*෎a�4u�4dT��#Ъ8k$R�d���Q�:���͉ϲ�"��$����r`�_�+�de�D13BSi��Ya߆�M�~�cF"V��]a(���0��xz�f�	<R��p�p1�L�v�[�#,�Eb�ħ5����Խ�<�P�CZ�O��q��� �F`�DY] �����,P�1I��_��wP5�J9`�-~44����zxJ׿��VH�`K��4$Y����]��5>��3J���:��v��0@g�� v�V�`�������#\����zLq�|�w/U� >>2ӑ�`j�*��Fm�K��ɟ�M��l������L��L����r��	�}��b�������,b讁��n<�K����j���ݓ��]-�WN���zQ�2�[:��GH�z(n˵���8c��N3�c�+=��V3̹����\ �4*v�u}�CUy0�eJ#[��C;5�@"*���(}�q�3D"�m ��Kkd�bT1��x�%�����2l��)�)P	�s~�ڡ�:I���`mx�0:�`��IX-��@�MھjR�������DĖ����5��RL���ì]�}"��5 �1	��j����p��Iw��W�Xe�)�nU��YYA]UN��_�3hZ]w���(�!�%@3�3�=A����"	�E5���f�������=Cb��{��%�M~�1q�=�T�S+�~�֗h�������������d:�]	�����L\����n��R��7@іZ���Q���A��N@-�����!�=�\>d�[�?2@{���ڶ�DeV��"5٫W�F��^�o���3�&:����û�>u+�7�ɣP�M�M����(uz����DVy���:�%��x*��O��N�#V�5*Q�e2��谖�S̸�vQ�1�ѨS�9�f��\��i����_���.�F:�c�����O���zivm��_����p��6�P~���yy��g��pR���K}٘�b��]̭ v�W
.���={�r�Bb���.V�ܴI
����Î��,�
�/uE�J�<!�Ơ2|�&�K 1h������ؗǦT�E��
ᛞB�����'��X�0��WxcZ�8d���D*%�K��0z`�d�=G`���.~~Tɺ��=��,w`�\��iS�5��p�e_�����5�W��&)oT��������L�c��uӣ,7.G�����(�/�I���K�H�3�4���ȻH���*���$����M�iXHYo�b�����H#Cf���*a�?�2{�t�w����f�PL�V~���śD�A�mN[>��"r-/�*qq�l3���ȝ�C,�g�t���^e�S�n�R�� г��(���Hvq�+�ۺ#������O�sb4GG��c>��B�砥zE��Fh�#�&���ݥOp��#)�Q�'&�]�Z�1�ϭ����M:|���#��w0�m'��k�[Y���D~b�aZ	L���򵨘vqR$좺m%dI��9o�iv�
C6�6? k��z�i�*�	|0=��ޕ��; �0��T��\�ի�V���\��5a&g(�ɱjS������)���^S�?�K>���٧����L��з��8�ٌ��KY[Mp<a�d����nb��
f�~�;yٚW]��_Du͈	'J� g�� �8iWo�Y�Lƕ^w�^b�wa+�� H�Q����O�����/u��:M�oF�ߕ�A)c%�r�Z�j䁥^>\��z��B��.f]��h/3t�/�֪u�N`l�p��'IMQxL<��I��3%&�79@����OR��ӋӍ:%L���md3!��a��&�]*顬�qʀ5�nqX 33^��	������=V$��~1�f��3��z�T����z9�G6+$״z��^�����;�*�l\ao�l�7���b�%��P��}�����UL���n���D�LMgry.��o�l�u��B(���KbdpE��JWtpb�u��tL��^ #�fӓ*���j�˾��sa0G�������<��`w�V�n�!4�L4񵘼�{���8��{t֒\NFMK�n��.��o� ���(Vܙ�64�!ڸ�$߬�������7aai��[9�C��.*��t�4ݬ	��������`��.Q���	Y��7)8hv��î�]����:��~4����a`ʬ�4��0$LB�2-���f��4:�o�������F�}?͖U&ta���Yن5O��'� rA�[�M^� �����=�]�Լ81�2�}\���PG<�>)������0Zf��8���
`��@���h�!���>���A�`?Щĥ����%����tHv�
p�/��2j��/�6��"�TͿ���܀ ��`gҺ'�$�����%��6�T�'���r��!&���P%2D��c���m����p)�F��o6ø��p����SW\nP�+]G&��F�ث��SO&�g��޶Jp�L0��=\6�8e�.o�ˈZl&�� [�u_ʍ��Y��֧&����r~���+Tb�(Ҩ��0���P�����U��U}q�r�Ygm{Ʈ�_K�ԡ���0t=r.�}�D��,Q� �1`<�6f�{oT�ާ��1X_��mQ������"�;�`���Q�>�׉(eOt �A�M��/����I�	SlA��a���0�z9(?�%+���l34S��xI���1
��2��n7P���D��p���$�xr����"��砹�x������"$-�Hd�v�a�K\,�x&P�}�")�Pݜ�Q��T.M����w̮�g�@�g���]���qy�!�Ls�9�@�ևe_�{�~�wQ��3���8ln�1��=���&��~����xk2q�:42P���*8�v��>���ۮsnide�Y~=����6/���S/��P��Nfb���YT�5LWs�`�����<v�UP-}�c����6��{���b}�3�y��}Sd�;��6͕Lp`dܫ����n���d���ܑ��_NV�{��ǡ���iը�c���tZ̺gW���Y�->������U7������$�P�a/�S뺝=�z�M��φ�e-�./��{�u��NB�Y�y���FE7R��OxU�2�?�G�C^� ��X-`� StN��20~�c�sΛJ���_�5^L��đ������3�y�X��[��-�Gc$:3��vڕ��w�G���C�G��YAEA�8O��*'s��%����b��y(et��xaD�Y����;
�ѡ,-���2�K���[
�nEpBz�����G�&��뎄qz"YA��Uʑ>�j���[�Y&(�GF!ԝ�{��~�Hw�y�"�3��8�n��0��f��&���+�ru�%���?j	聶2( ��ۧ|) 7�K}7�}i4������O�n��H�R>s���w)/�iۮs��Ϙcw�S��L؞��!�-�AK�c����qnY9��\�hn�-�կ�%g0͎�ci	+�v�x��("����)���=M�}��l\}��Kk�9.O��(�j��r2k1r�.Y��DVЖԬ�u'}��z�Y��]$��:�Ѳt���_@O���Fq�.^�>�4�iY.����Y-5��=�0�%�e��K���V�I��<\K���_�~�h�A�(�P��Mb�)8Yt��qsa��^�?jF�hrΉ���Q����ˊ�3�3L?Hjn�����R~~jeUJ�B�ݽ��է�8�@^��I.��V*o�	�`�W]��VT��֟��-�41����J��Q��i���;�M+Ą�R�N�@n�2�Fk.�6�
0��p0�\�,��-O��n&��oj��u�[�y:Am��F� �Ѳ61�,p`,�h!2	�C�`*�)݃�<KP���](��\��VҌ�Okb+�U��hwr��3���J�B�kA;�V@ ��]XX���5o/���q���$}�?ɘ>Ct�3��y�R�wt^��A�������9@��������mQ��a��(����/gsL�77��^���c&�Y"R q+�%@a�eǔF�v2Τ�^�Rp�%Ւ��Z�uHy6נE�p�Yu5�"JB�\��S
u���A���I'j�����2�	˦p�pچS��h�"�:�2� ����H�
� �ti����L�4V���� �G�(AB�r�Q��9+d��דyd�u�4���Oۦn,���9�.ş����V����(�6���I��#���|m�g˩��[:�UAM��x��h
?���H<)�~������G͗�< 5x���ִ��Ǝ.�����'�ȓ-��c;�*D�	*km~�t�1�<�0ʆ�G�4pW)I�X5��'�:S9D@�7C���|�N�⢨�n�s-RZh2t����[Ng��_;��J���N4.�G����~;~�I�t\S���������r$,�:�W�v݌�r��>�xT1��t�J#����%��y]0�dt.Ǹ�y�����n\l���~P�H����_��I�`�B�,Q���?��͑X��$d�ق%��éf��(0�̞�>�(����������J"����H�nP���Z���Q-���a�0�#�Ƙ��C�Ll�+y���>w�a��(_�j�oLA*&<<b������)t~Q���z��U�q����胄Z�D��k۫R���+�r�=�i&Ґ����vn�.�ڦtZ����q�+z7aſɈ$�i� ���L�E�h���,���߽�vr���n�%AE���=�.�`����cR3�*��i.�wR��UQ�rJ�@���n�nq`���0����.��+j�-0�w�4�jx��/�ld�xT}r�,R��w�]\�G�ӷ!���gH�Qi��0�7���L��[�p�'CLhs%_�:�?��d�-���e=�Q(Qm��@]n���%YG���n(�o��y�<�lЫL�J+[j���W�p��(����c����j�
 ��O��0F���K�C��� �=�����{�DIZ5��e��9�߸I��RPD��-��&��B,�*R�Y;�\��!y�g�/>ƨ���c�
��!$ı/mޢ,9������%0s�r~d*Y�s̞�l���}�!zTMR*��H�,QMCK%�q��IJg�2�rE!�˶�1rwx(�\��I! �؜��G{Vx"e'>�/{.#r����]�Y��)���3Ku�5.o�^��q�%�<�y��-&�e�~W����q����ET�t�qE5��}vr�kf��|�pPv��g��UPAɇv[u���>�&����U=Dƕ�C���w���Q۰]�f�}R�z�ҳ�2��y�b
+e&�k0� �T�q(8<�8#XT��_H�u��>Jme���H~��د?H�A�ee]%�_�Y�Y"�B"<�����I���8�;���t�8׌�-���ږ�6<�3n���������\��6s�/��#���Ԗ�������\;*Dx��[�O��?9w�tj舜yK�:(!�)���/�[bդ���(������l�ҡ�kp�ͭ�Z�uH�ĻԆ��V~����Y�����&Ϋ�ᒋ������Xs.�q���*����S��&Ƒ��q��-Y�}d~�G�R�C�s7<fJ�Y��Dʥk�0�9��Q�sܥs��,X��ET7�W�%@?��������o��_��ɡ�_�g�8��`�	�ӿ��x�����x���� OF�������-}.o�1�8K��`&�} 4!OBu=��2sڰ�t'�����~��6T{-��mAA"�����p+�8^�߲$���I|,$��\�#�N�>+�1?E*A�}��?����#�v����� �;�y�"r�[E��/�o�����@�2�"q!�o:".ț7dz�V��� Oؔ�*H��&��Aޤ�v){t�S� �i$����v���i��L�����ҾqfS�XS�6�H�t\�J�Yxa�O�/���	L]:g׀��=�)��n�� �e�\m��B�P���"���l���
����,�DF�s�,P$[l*�zG���r`K���ݬ���b�"E�l�V5�CU�󗡬�QBxB;S(�/Ve]�^��@��7ϗ���W�u�!UA|���"p�+lr��
�x��t��Zb�DtL
iſ�F��m���o"��[���tͼ�{L׀$RM]��:?��"���]�k=�tX����I�Y&�a�� �`��a2��b2�p	@�{z|7d:�$��Zb��/�j�U3�;��K��o�� H�N�9J�p{F��^ħ[�~��u�~Cm.kA#�I���vJ����Ǿ�8|?���M=�0I����\�j,�l�7��D�N���9��,�a>cT���"���af��[^s?fa�Nڇ�������u�y 3��Z��ɂq��b&��vc}�>7��=���@��^�:f�u�6�����0!Ɂ^�:>����� �e�n��ȢI<WS�9�p���N�(p��i Zϧ��C�'�| �i:�����\��|��,�}�����E� 3��tKvՄE��;��'Uu����S$ &#/�k���S)p�]Iܺi�"�[$�Ч>�X�H�]�
P��!Z��7�Y+Û�m�=>�M|��J�搔�~�Y<���VBO'q`��Ѡ^�??))?ᦈ����4�:8ʏ�D��{�~<�6�\��?dԣ#�I���:;�6f�j�GU,2��u*����D�&O`�e���F&,j'���fP�lrv��mQ���}.��X�J'�������j���g#<dC���,7�g�*��:��Q�}�B���5�J~��|����Ț��g-m�N4`��P��-)�֔�6��!�Թ���Xd����S���ŏ �-$�9y�z}��l.�	b2R<_~�$e/o�/E|\��~��LLn���J��#�T���cA6`������Y���W�C$c�g�H9L1��{7�ua��<d�+�A�7��p�Ub�v��]h����/9& dsL:��V�_hZ7�����6)P}En�Ds@��t:�>���qNw �p����$� z���$5�k�{��ϲ���)�5 �i��d�Q���D�X�@����P̆#��˶����YV\/li�w���~NK���F��q�,/���j�m��.FQ��Z��n7���s��O�d57��3�u��NC�؞j�0D�-UcbytQ|`b5zP3�5����ka)�H���D���L��)��w�� ;M�F5�Be>8F�㜱s�Z�J�چ��:��CK�I/�>�$�g0G�f��'̢�MT�0�^j��ɦuj� ����q�35F��=�Ӭ�(��!�?��-��(Gt�F��Y(4Moǐ�������#��ހ3��J�S��Ϥj1Cju�^��{���ވ�g�r�w��"�5w{9��h?���]DE	'�5&�@Ǧ\e��_|
��T����	�sY5}�3��e?�iN>�iO٢ 7��'(K�-(�D0kU�E���j	]H�P���u�4�si~x�[_�l(`�C_�Z�d�H���q`fR꾁��Rp���)�Wo�i��c0yq���L��%rA>׸�*K�*C�������>,�]4~�^��-Z #���%�S�^��ŕ-XlxV64EB    fa00    2a80,Z�begPhv�I`n��$B|��γ����;�u���=��,4��"��J��C����	���@���y"祈�S�{XR�GrP�9V�z�_F��!Pw�3��pr��O�=��������"+�����K�:հ��sSh|�e:t%�8E]���C%�G�K�щ�%Ӗ#�I[�9�W�AB����q�ix,6�w*1|?�k��[�A$6Z���k��pJ�Q[��A�8��$�GcU�����߆R�D��a'u
���?c��7�o��ݶ�;���Ao������Х�������}�`��G�������2;��^7@��)���K3�����ߦ8��u�"�1u�s��@�A��q�##+� ���K1�A{����(���D-�� ���g+�G��<|S���"{v���ȫ��=_!2�Su��g����c���RãȮ�yF\��;�'���w݌]�
B�K󐛂���1C����^��\'�"zJ;�P��4��9����o��`BA��"�ۉ2��h�9�|��PB�w[�0��(��4�Eg~�Μ�/b�ԺK��7h��oW{Q�a�U�} ��Q�^v#K�;K�
nWB��V���b`O�z�Ek}�������Se1�����\�LN�D�
A��'FՓ�f�-��$&%�,��_	ʘ�z�x�E;��M��5?��8�$�;~x�x�DJN�i>BJ(��F)��)���-�����$��P	kֿ~f�����D�5����d�����(�Kg)�\������>���5P�����b���Ly�+�. ����
RB�v���<����w�|H� a��o}��Rm���+�����2��bۧ��[!�ws]�Лb7���d��|���ێA�H��u<�$����b��k��1���F(wsy�S����'~�ū��3[�z����#�>)��8߷9��\�*�����{�vi48]8�2�5���w���ʃ���7:	5s�;���ՑC!�;�R0_��ל��3�O����!����0��ÈM�����1�^%��qM;�dp��C�-���0&���P���ؾ���{�$�L�Q*Q;�Gh@ɪ��O�<�f��-����E�6*N%�������qJn�4(m�:�&:��s��s�H��٥��9k���'lre��P}]�ke�(�l���U#���Ö_ q��D�B��!�g�K�}^�����ś���"���J��mC*�4�Q�m���H��-�"�I�&t�G�-z�oC��U�4�Ǐ���>	L$��Ԉ.W�֘�t%(�~s�C_���U/)��T�2�[�v�ەe�>4ܠ�	�{/��T��-Q�0֮��z��͟�k�z`���ɛ��S�UB��������J���9̬
�6����r������s�C9h�$	唕���5Nk}t���H��m)r�����a�ٲ�㥎1Ĳ1�ʏs�m4;?so**s0�i&ԟ�ɼ�����T�Y
���W$dq��em� ������d���7��(O)`E0@냅(i �yհ���2��#J�M�5w�n��<�_L�������~}L�+��^0��*�m��{�_hP��{���ީ��X�Gf��d����Cf+���bDHlL}��~�J?�Bz|[Cƞ��d��/A�@K���،[ڮqEW�{�k��
_S���v��ًd�v��2l"!�uǌ�y�[	=I�r7F��=�L�6x2������^�H���ا�P^S�مW�S�L��,�WiyZl$����q�}jj����d^���c��(e`8o����`'?�^+\�vl�)�,j�B[2�'Z�KDv������'К)Goy	��̈n��~H�(5�Fb���w��5B�Y�f��eD��E�Cb!�㘅�#ڭ[c���\�JH�Ifw�Lic���@M3v@�)A�����O�P�a���i�� �8� O��D����-��2�Y��Ct�}^��ѫ]P/�߻ʡ[2H�gOx�H�HU�%p)�q�^z8ePj~BS,���E��&����5��fX�|���S��l�E�5����j��7ͬ��Q����t��5��S����d��Ɨ6s�˨�z*Cm.[�_Q��.�����S ��-rx$*sFʻ��C`Y��4�iiIؚ��3�Յl���!�Dz/�
��j_�r�K��c�'d1^ S��@�����\�bx�����(�O_zOP|��W=����x��>N� �^յW���BG�A�u������H% �7�l<�����8��m�J���VG��&�\N&*��8�Q�0�6�����oyJ�[6�)����U����Nʓ��o�ࡥ��ƨ���cx"κ-�԰�ֲ���Х�\�1�w�	�|��.�Lr��J\6ូ�I�=B�'~�K�pR_w3�Dr'�u�hE�x8���9:�sT ������">�sb�5���$���J%�2:O�!#{�<�,��VL�E�8XL�[��y[r>@�q�%k�1PA	�x%���B&���t
�Z⊵Y�ϊ���n��7_r>Q�{����F&"8v�(SB�P ��}�;_;h�]���p띓N���T�DJ��{l�eO���?p ��=u^pq#؋����I�,�t������ � �2� ���NC�CP�F�(貚T��oO1�kc��_!���r�|�]S
%Ă��SD%��~`����WP�Z`��&�1�9��R����|W���iX""	���V�CZ�T�u�P5"m��/���\%��E��	@<n��G݁���Ii*1F��/[NR����G�Do`NI="\#����'J8_j�]���Df]ң��d��rFTY{H��y»�dϭK���o�"�υ��1196׾O�kd��y�T������<Nd#B�{��ra��7���5�h����k�w9 ����z��l��:8�E��7w�lcT@�O.ջ�Fs�B��	X��z��c��ђjq&?���~$Hkd'-

��O��z��l!X���K����=D�!������J�q���v�M_��=GJo��4l��Y��.�*N6��6C��^���%c�2���/+8K�.��G����9�ѐ`��p��B�ʓ ��T��Y��αIF�]�ť�ܴ�9�$�CK% t&�Įi��*3����8�ЍG�(%Of,�J�ţ|��4T�9Zt9ԕ���r>>J%
����M���~��<��Q�ψ�",�?e����׽�C��/���gR��	2 ���2Z)!:8�c�����q��㬯D��ՇPI%xZ�r}�������)�09�Fv:�|5~L��u��۪py�o�����[���|�Bi��'�6�Ϗ�t�M�ܗ�r��9��0�VR�����ku�В�]��s$|�2m��WT�]�f/�1̚���@�k'(FZ�<� LG$M����Q&�J��qpC�Ta�uD�e��2/�M܉��KȮ��}��˰L��N4��L@�ǊL�����S/���w[t�2$�Dj���ĕ��3J N��\-n�C2%����Ս?��(ʹ�-t�Y�u~�a.� a�E�%��XI��(u��W����(_�z���C"˛��� :�&�=�r;��V�4�ڍ�C��}:�;BK�S�����e�s�6�$ �͠��V�D��"��Lnz�cd4�ga,UF��jS��+T3$����%<zf���di��@�	;�'�Ex��A��q�Y6�����#�T<6_�tF��e�T��C-���2A�,T�G�3�#���NI�3=qu������"s�_m3��k�9+����zL=�e:�8@0�p=�\:�BE�B,�,��ꊀeGL����o�5Nѻ��2�RӺ��l#���a�F�3�/���zI4C�߉VFRxkA�n����;�̺���,H��T3���M5���Q�uj�>�T��v-ҏc��#~����
4q���Q�鲌{������ס+w�%������m@5��$�uc-=��ȑ�n�Z;��@����7=�|:��8�l�����	��b底�n��A�ehH_+���7�2k�T���КEY�$�$�V����z���\�1M���W3קy�V!�l�+��2��Ɲɽ�!2X���3o'��n�ӥv�}DB>-T�xh$�d�+�^�Wu�7���;YQu#$�+��.k�Q�~�@���1����'�ھ)��~���@�νLy�����ި��Zܐ9���:y��I7<���
���r}��ͳ|���V��������+�]e%�-��?=ܼY���oP�̀|���%'��nD]����iO u���'��	�f�&�c|�d�RV]���#z��>&)��	wTa˖�]��x�>����(�w�Hiϑ����VsCD�s�>3N��T��wC3��|rN���,j�:�~��X�lG���%P��``k��,X�5�ߓ![�t��@5���)�
�!�|��fզ�,vB	=ү����}伶�=z��L��J��t(�����x&ɂ�3tY?ݮ�6��j<9,k��x�n.�N��f��X#�H}v1����R'�,�rS��03�{�6\/[�*�d���J��`Ȉ>��(���A^zsǢx��TtBMAߵm��|\~��i�,!N!��<w��`vMnQl�����o|�R֭�f70��w0�*���kS�4��	���0�i��2hU[�����#i,��~���M�6&vs�<�����n�Q�/z�^x��SٗA�Ug��hw5A���\Ǜx�d�!g�K������*���"�c�D�2^��R�Q�V��D{ɣ~���������s�e��BCbfЈr�X9�9�M?�_�=��ٺ�#�R���,�4W���Xt7�|es�d8��jR�.�1�Y�[S�#}��>h���������z�J�VLIev�Q���R¿�Uo���r�f6ہⳠ��5*M^Q��u�**�x���`��I���X'*k5y �:v'g� A}a�ϓ���!��U�+F�d�4�d+�Xa|��Z�>�:����ǒVd��u����O��'w�XqIE��e[E�xv�E���d-�`uL$�2e�#��d��\�3�U��T�"`v3�c�Ad5�$w���R��f���5�}��J��F�AV�5�Py�G��ƿr�����;�UP�S
;EFv*�ǌl�ǎA���n�X�Z��i#�nѲ��2w}�U�f�~�3!-�̜␪��GB�bf��8�������JHeł���:���"�S���ǊVU���K���q]��dP����NXN��M�%b�Q���L_N�
���M⬩�T-{6V�L�;N�r�mse����C����i�c���x���7.?�K/�~LQ�&��FZH��V��A��
(�p�ɳu8�6����"�K4�&��*���5׈�� 
o�* ;}��+U���q�Bbz��ivȉ��*���cY��Y�T�$d���Z��<{�Ģt�
Y򨩈4N^��C�.��Ht�̹�%r#yuj�c��F� [Wa�$׆6]��o_[���������=٧�3�Vj�&�AD�L/x�m�*�����by=`)<����N�;����5l�KLB#��`c�	���M$f�.����Z�P��'_�;	��J�;}��)��7��y���ˌ�����A0�\r����B�=S!ӆu�C{������9cB�5����WJ�l��|�W�m����]�?���@ ��1��Jp�eݘ@�I,����t4��l��%���?���C��ִrE3��p�X���+Q�2�G�3{_�x?,yAۼ|m�"���=y4�I}=�� ��^���Ň���^�����ɨ��&��8P����/3V�/׿�>����~��<h��4M^�z0�镆"JƝrfBbR}�W�'&����0�E��Q���5�[p�۫IՄ:��|>i���(jcG��u�1�����U�G�q�QD�;����P����CǔF�^Z�~ŝ�	����!$Rr��9i52Z���U�u"�q����9�\�YK	&���.*�o�1���Q��:)�ԭ��{ۻ��.66b�
iV���-o���1:���I��>@j�;緘����M�$މ����D�)^`�/
ſK�R��� �-\�9>(b�mk2��Fe�SU��$~&[Q�0ޜ�fL0XM��{>���B-po5�Σ�B߭��(��e���T��P��O*Q�'��(-�^>Z����s�w:�O��a�bw#2���(~���ph+�s�9�*YdKQS1��&}�h�/4�J�n#�v��$l��	^$ȽƲ��u��pZ3
��������_l#y
M�[!XƤ��nU(�z�~-�t~'VU��L
�:�}y�&�e���-��_|�4���g�|Pa�t�E�'����n���ϼ��t ��1Y2ή��Zfʹ*w�_�<�H��T$C���������K����=mr��t�7l���	4נ�"���<����X��Z�j����h��yu��&Rf%�Vl7�e��b����K�[u[�W�Qz)��9�8"�Ԭ���K�>�,J��#v���{�����<qNid���n�:xj4T�A0�yӆ�:z��h^�h�H��%�sky�̅�-���9����/���:!Byډr�g�����+�'�9�_�tMne<������j�X�^W܂�|���3Z�����l��t�v��9�x�e����\u�f��qx�WcR	� ���A�\��&y�"�K:h�.�����jLל�g' ΐ,Ҫ& ��/�=�X{�u�ȖH˅L���bH���E>�}��i������/q��_yNvv�A<ց��\�@98k�ū���j����'�, b���<���s*�I��{(�&]+��|� �'�kF��]��c��7�n������!��>��9��l�>M��wu��(�Q�"���j����=y�j 
[�q�KD��=�k�ib��bZW�XÀ��zL,X���m����'����!���(E6����'�k{�~��a5�-W(��3׀[��V����[yA�׮�"φ��/X�7���^<&Ğ�
=��|�b���*ܶYG�
_�{��C���!����?��SN
�Ov����K��Z9t<��#�X)`'�m�Ee�<3��h�PY8s~WR�멂CÃ���E���ue�ƒN����rXu���Iqtɩ�� ��Y�	�'��=��R��d?���5.C\7�ܬ|�ӿ+xF-�9OЎ}�.~ �Ô�IY,lH��e[����:,,��J��1����j�F!�<�$А��CA16P�x��!��/�.���`�c,��*����!�Q�k{����p�r�h��^<�(��d�[��R�RU�5���U����T�)�~��'�����܊�SO��C�� a<e��F��{��F��HBj�#)e��7�K�����@��J�j,�]H;��Tg��r���~�xˆ'3%8ğ�C8���� z�.�ᄽ��*Ή�����O˃���3d"�"����8��r�$y���[�AںTj�8~p��l�ٕ���x:0Q*�d.��Q��.e��ƯZ�aL&��UP�d����!u0��{�=U%�+)�
�Pa,�J���R o΅�9�R�R�oe�9�m1l��V����A�-�������y9w+�{��v��;����;R��c�x8�
A}l�_xǄS`�2��m��qJN�v���U��b=P�^��{46ކ���6�\^�2;�����'�3:�C5<�	�ާ�&WQ�WNR�q�D}F�#�{9���n""������}#��BцK�^J#�Ǖ������~��X ��!����Y�X�K�{�0���i�(�j)XM+�#�xB�f�K���8�O��KP��FŦr�`��W� ����)7[_͇��=M���a�������gv�Q���Yu��d:��Ҧ�0w$���uy���S�
f&J`��!�&�O��a��>U��t�1��-�0hK�B����A5(c�G�7\S8���B	ie遤�Za�M,Kk�������B�J��'�vm&QO����F�Y(%��K-L�0�1/��\��a+��=�1׊�N��E��ު�u�u�1%/rJ�c�
�UPj}��%R�E�+�r&J<����a	��[��4��х���o�&�WwȞ\cy��z
da���`���������0�Ƃ��C(r*��"�.���=��:Q.x�N�	���5�	����B�\���A�>����)��[�`�u��X�"D����S3x'�����t�v��_���&搤>y� )��^�*šݨ
\�� %���2#O��c��{�z����I���$�ÑgRP���K*h�^<�Y}�p]�����O�����D�'��l�ڢ�>P|�MP�I'A�K�G" ����ǌ�8w�����l���!HS��2�Is\kr:In���|_T�Ӷi}�ަ�c)�1]��A?�{寘G��J$l�n�O����	څR��'��`s?����l��A���Ⱦ�k���b�#�Lt�����̢�kA!�o��U�:��ah��P�p�8HY$�F1u�T0ث#�U���
�F��U#�z�`�R�[Zۓ�i�)��z�P���3��Y�ol(��9��}�e�90����F¡�D�������=���i̙	b��o�(7h[�����OJl��1[@��r.� #�������̿�eG���1f�3�|ؓ����Lګ-M���7r�k�����v�=��ls˯�eC�%�M�m�όV�6S�Q�g�!|m['cʬg�����ް��pinR3%�L��+ �y��ݒ��s9��(�9(�S�8�YU�E�X}�$e���NG�0����˿��3Mc�\lm��$�gn���?+�i���Ӻ7��7:IR�ic��V��eV.�H~:Kt\�q]�;k@A�^�F�xXK�I�3��
�������K��gY����pM�d�ތ�'�^���8ٿ-���E�"9:
H
�]�ٲ�1f��BZm�R	�=x�k���5�lW�	�I� �z;0�� [�����51��;���熗�9�N;'�g�F:|5w�D!3�b���;�L�
)�Ub�P�����W�EV���H~Y�B䲐&a}�����=�$ӵJ$؏����`��@�K������y�K�ap�6!��Z+q�}�#��࠼���T�W�B�ǟ�"]�Cx+t��P_�v��n`_��x���ʦ?x����W6�jT�W�:�s���	��9�������x�B�Ւ"���9>P�
�O�μ"9�G�lu�xg�z7��q�Hdim�r&��l�Xv�L�o}�F�i�``�'�v�&5�
��#Lj��w��=̅͐��(I��[Ȍ|��P�_8M��W6�m�Q���3��: ��� �����K��qչ�E�X���u@3��<��#�]� ���T��df�?Ռ4��e�C��ſ�+�0���h��Hŀ��;=�>�$|�q�qo��ꟷȲ���C�Z�9C�%�r��m7�cd"SKb�\YG�]��}ح�x������Y��R�r����A�1Z�CI��h ��'���vYC���؀y#�@���2��A�������1��m�5�����X7s}?�h�u�O��n��'*Kz�|�@��O��s�$AJ��Gr��C�X(a�2U27��N֠*4i�(�pǒwǊ�
�-t��fGy��^N��J�́.���gL�<�r�5���e��Kk�)B��D�eO7�:�,:4ki�%W��2M`�'����0���.Z,)ty�����_�ǘ��~/����P��s�.�y¸stƤ���-�x�K�+�m!�%؎��F�YC�ǘ)�6ߑI9��!�V�v�s�x��Z�
�2��W��'h	�\W���lu�'T,�(��x}j�R�p)V�.���}�w�u��Ƃ�L�bT�F�僀���w@���C��IȷS򄯼����iM1�a�N���F��.���u
��DP����|��k[��ȵ4*��Z�/����i�NC�Ջ�24�H�HG��8�N�)Z�E �/�T� t`�$�\"���[?���+?k��V�b.
�G�^V5�T��h`�6_�k~�F/&*����T�7:d\faK_�����kfw t���z��%:}�|�Y?���5�&�X��������S<��[3�85>i�[0e|L|���~�4ZT�9L�J�W��Ge� 5�/G�I��)�S����� }�7&�2C��g�����BJ	�~�J��p/��T,ud1�Id�`p:��{�4e�b���5�S�ߔa|D�|�a'a�}8��Q�fB�����ᰠI�*�(��~o)��RFu�wj���.��b��dT����ȵ`��wa,�}�
��9+����	$���+;� �+P^\G������+�A�w����V�}�dO��6r�ZK����ۡ!j���M�:��Ba�a�">�*h�F��Ii׭���	�H7`��*�Pܛ뉻�.20���`��Q��V��heb�e~h� �Z�ɒ�����h:���頿)�XlxV64EB    fa00    2b80�H�)Xnj�A3û`R	��M�3���h�H��'��W	��|�\�r�Z�N�͐uqmǗ�,<[̕�m���[ԁ�y�D��*tq=7��3<�yI�ӆ
���}QC��Bf��_�����X�X$�������s��24��j���ЕQO�� �<��ڃ�)����^��<�,_��=\��a�ݿ>L����y�ަZ[����^ق�O�7O9�����-wmh���QIQ���9����K�2��m!�,]W�k�ѱ]�
�9��Y��֊��DeW��7�!a�5����J���^��V4��s���;�8����P��*J-{J�Hv럤�L@�U�,�5Hڢ��<n�~�Yc�csmc�$QK�����w@x~� 7i"+��������vH:OR�|�p��b��N������6��TQb*6e.�y[+\Z��xə'�w�`O����g��p{�I��,���IEw;G�����3�(���g���HA��έ��]�x9��\��#WL��=!���{ �\ϺHl�n��[���m��f�a� }�lk?�k�XlP0���<�=���*����7l�����|6���)V�b������ y&�;�~��\�8�J���}H%���	�;�6\��ÿ�NP��<�D�6����D�E<�O��"��6����튨�P�թ��Ҡߠ����X�B���O��d�^AA��NFв�(m#��ř�a8a����4�4N˃_i"�}���
�:tT��H�sg�G+0x]Q?��rv ��F�g�}��v��g�m�^Tد�ʿ�7�Z�]�t���=*�P��x*]jy+���V��\j�d���Y�tOG�p�f7�x\���sTex b�l/�L�r��U�
����`���"���DQm+ �e$ɳ:��$����u2�s�W�z��Z7s��94�ȥX%��T��p_Mx�N�O�.;JN�{��$^v���|�8�0/��7n��y���"­�v��ݏ����4:mP=���nd����,(9�i�GJ瑶5��4u� ѹ_aGN7)"�T=�H2Om|�a�E��������"���z*�ٙ��T�W�F�'(���&��{$��+>x
���k>"0ld״(�}L/�E�{7����Q�3I�)����d� ���DJf�e1u��W��4�S��q6G�Hx�vX�\{�nJa�{���?7�d��%���ZT��h����ij�����q�tf5L�jt�){T�
�8���<����3#�_\'<V{{8�*�p�`������<]*y���ԏ�~��>l�k��7�7.$�`с�D=��ip߿\���g˦����7�v�g(<��E��Zf�$�*ҟ�/��(�l���E��~��Ɗ�}+��0��u׼N��8�"�Pii%x�S^�%���͊/�R	/���I��>�eh6�ߔ
х��!�"�Xʹ�4��df��M\5�V��,͖fr;�P7�CE�%�;���l ۭ{�d8C�����;t-Nwi�DO�!=�%@�9�L3���E�u �� �㟀�C�t�yX��&��g�/���/Ύ��-�� ᨅ����/������;�6v�T��B��s�5S�n���[ 4t��B;
�8�q�r'm��� �}ۨ��x��A�?�x��ǘh^K�ݞr���j�����=�)��(�����&�]����,v�|�S>#��&BS�J�&��+@�Lo��?#U���z֕!�Ŗ5ן��
�$�ZƏ�?��[�ї)�b�i�!�R7't� wN%���E^o��q�2����(�Fڀ��^��T�!��;�'��:��wX��yV�T��f�z�<V����:��t�@��b���+��
7�_�S���� �E{~	�����u�I���`����c˪�������A�OT��8,��T�`0Rٚ�E�?��Έ�!����9z�F_Ʊg�^�2�F��7�N�簶"�<�	˰8P7��P���X�����-p'�6�b�ɡԊ$]���^�X~(�sMS��b���(#�"�����,�*}��[�	VC�F:��	�z��a�i"˟L�ȐJ
^��m<'e��ZD���� 69�'f�����uoM-�?go@q��#NY��H�~�ѧ�`s��TV�Š����*���*/�/�[F;e���x��wm��厼�f,��8l#�R�փ�5����~z���\�Ϝ��B��TJ���C=�8�/�np���,�n|6eN*2�O�L���$_��m}���p�|P�m�1��$���p�N�,�.A}<�� B��W��]PnY/��X�����d�LK99��S;�����9�G9��g4��ɴ�H�C��;c7�� �~
�wo%�,e~�ɠM)\H�o���e�囪X�կX�{�8N�7��Y9
h����U������m���M�dF�~ �HU���>05�s�t�8h� &�*J��}�knv�͞��V-Ő��'��h}��F�b����O�~�z�Sh���2O��9/�[ ��(̷4����+�d�,G1A����G�H�_���"d��R��b}��>W���0mv�2���.י�-��E�����/��k`"+���oR���5���N��F��70�e:���V�s��mvԽ�2���*ZL(�D=��SD&��-~]_]��E��P���0����\���v��%xqa'���w���v]Hz��~�/���
�_�A\�/<��`X �~���,z��[���WN΅hٟ�N����Щ�����l~BHg��n\�����@��u�C�B`�NX2˫�9aXx�f`P[H�����)�H���H��J^��R�.0&2z]�~���g0p�q�	b�1�-����)?�ň.8@��Q�������m����P'ղM",��1�g�}uG�^� �^�����c1��	�X*h@��;�&�7'O䀻|�3lρ�e�[0Aw�-ND�2��D���9g�`��)�L�0.I`W��H?�D�:��\���������{���q���`�o �m�m�Ec��f�#�$WK�A���[�5��r�e�;˚�!�3�����G�x5�����4&�T%�����է�`�ǔ��$�E�p�ta��O�{��^ʶWğ%�E<]�a��p��;7s�0MX�jJ_�n-�y�Cz�\��T�LT�"O&�YJ���L�JY
"���w�94�?ТN3���|�ӄ���@~�����aip����)Yh���4�+�E��i�IJ9�7"��M��JK�-H��H4��t����"I�����9�۴Z	V%h��|o(�]+�B�ݽ����KFK�,2��	8��~� �U���g'�a�bY����QZ�I����/u��xJA @X����E���+�}7��;�c�ԯd�[����~�V����q}_�=Y`��{Gc1^�s����B:���0��\1����(�R�ږ�-�̸�=]b� �1X�Ԕ�;�D�Ϻ���/8��D��J��J��*���!�2"�D�b������}�3;6�yZ�?�bhɱ�s����:2a-���ʋD)����Eچ��)2m��d��9-K�c,"{H���<�C %����ƚ<ʋ���[<P����\e��==��\���źi}2�Ҙ�6%�eǝ��� o�,��2���9Ҳ�X��rQ�������>}�����IZ�q��C�L��z�vE+=$v�{�hfe���\�ljQ�������, j��&$�j�`��H��9\X�X�T���y�;��i(�I<O?���R���
�
���c�=�{B�i|2�،�E��B.a�c���������0�i,��ؔ���Ni�����plr�N�	dvn��;P�%�0�u�]��A�6H-#S͹$��J�wi�dy�h�N�<A?�s���V���a�/��t�!�v��#�Ow�q��H���7��C�s%��+\���ɰ@�/�_?�0D���v���/�#�:�4T����娒��Ϡҙ�FG��O>��G[��Z�6H�;#��i�EUcbZ����	��F�
��௱p�P�D�y}�W�zDx�XB�r.8NQ_�7�!��,���w�"�(�$��#��$��;Z��W��6nj��cR�oP�L1Vz7�N8�]�����N
7M��#���ԇaA���>��9����l	��K?)�D�`���D/
|w��=ݟO�%�柌 dT~�8��ڇ����^�*,�d�
V�?�y�T��6w����ύ���il)N����4"�2):�AH���Y`=�ƅ -�����=�9���ޕV�2hSk����q���Am�t
�%O����� p�V�� q�AD"�}�����ȏ  a���1�@��@J���x@ိ�h��1�E��C������c����q!����,�)�"z���� ,R�BĖ%O[�V�?�`�<R��ʬ_�uE\��zn2���,�dfC�J�A5�Vσ�'�+]9᪵�(�7���R������b���bF���G�#vy���%M��� �C^!��=��Ț��
��X~�"ܒ���+ҷa�C�3� I	�<!?�k�IP�
ő�������{�D��B�ؠ��S�:&p:��M!��.�Q�s��QA*F�ώB�LA�>�20�v�Au�
'\���~�+��������R:�����د�m$���4gW�?^Es��9F��.�P�����j�-�a�#�*=��53mt:�+�/o����=8��H~�Q�^ ��c�y��i�������c4�]��3�����)���T�������U�;��A������*5x��Ӛ2�i�\B�����i�Yh&WO�����u�۝�PY� �)w���\���B�3zaT���%�[Љ�%�N��R�@#?m��EU?x3���U�`��V/%����X��A��$��wy�cu���E!�]�d�8��5��:L�WKa�*�tk�j����-)��;�a�g���d��	1 ��!��U�T��~���Cz��"L>��_�v����X��l0NO+�.-*�M�������
Ŋ{"����Һ�@��2r잁�@_V<<G����7y)���.^�r����
/'O
�\e����S���,а�n��DB���7�ƅ��o��c���Ǉ��pP8���D�F�6�f�֔fVL��n�Z� ��)Y_#��k��0b�sT�(G�.�#ņ��/�e�G��9D��,�q j;���`�2�$��͸�dF�/N�S��Z���/P�����P�=����E�4TE��Y-����yv���։A�v��Y��������������5���(W/���Æbm���*���Z�^�@�IJ���!?�!�ڎݶ.�_p縴���m�b����(�A ��죺�+BV�6 b���� �Q-��Ҡ~��ȼ�/"-�k���}"��$���QOԁ�:+���K��|c�x�hoY���n�9W$R'DuйԛV��q>bX&���"���R,s3�*���IY��K�}rq�7ݝx���ؑԐQ5'|' 1���h�eI��]�c/�Ŀ����������Ŀ�u��l�	yHsaF�ݫ�I:Eɣ�Ȏi�b+��B���p7�j#���r��O �8�x� �<��j#���_��k\�5�6?�u;��'��8B>It�	�-��n-��P�b�{��ό*F�Ы�>p�K�΀{�ޖ�|�h�X
2����6c��1t�a=���C]~�ͩ�`n@C�����x���6y��� �j>D�T!P�S����cu$$����ԲDO
���ṧ���i���t�ID��'� 4��<���KI歴̏�}��g%��KmB�ߍ,4[l���%�M.3IԠ�Acy�T�t+ʿ������/����×���e�.��Gq��A��1�{v[@�����l��nܻ�͉��A>!�5ԋQ���xtѱ�����tu��ԍ)�~��ub�Ø?���Y�d�	���%}��"�{}}��i��LL���ý�Tp�����`�.4k�ߎ&+��C}D8p�$�F���/�1z>z���.,]��_ �����k #�fб�T�F��㑎���@���*K�O���I#z�K�7<���	R}������	%jt�L��?�����M����jҨx!�B}�b��j��
�Oj읤7s���R���Q�y[�k� || ��3E���C� ܏���p�)#���@csES��teA(�~��mEң@�68�F�۪]�+�4�ߝ~�ne����Nſ�&���Bf�4�rp�6oOqV@�-y�>-���TC�X�c~zl-!Y���4��[�I���VU殇�H�z�B	F�p����I�ݼfP��t�ЋJ35F�7j:2�Z�.nB�7鴸>��swu2���"/�7��,Z�c�8�u_	_�������A�:`��@��qƓN�����&��G؅O���2������y���E�0&���G�%�(��q�S��"c�\���͚�۵�%���\U��E ˭�̷�.�8���*��-��*������&Ͻ#��9�@"	����-#��fv�/����@�u\ȫ�A�S����v���>@&PCwC'����m9F@k>-g�ӭ�6KӍ��Z����I�iJ[�mv��/2�`��������Q�i3$a�`�H�����D/:�+Lٖ�Q��,��3�YS���! �쌹e.���5Z�<!�s�3i[���~�@E���t���$�G�
���ݢ�C��
lc���UI�y�+ې��~�fӠg���Ss�|+˾�_��c�������q���ލk	(�ݢU�$r�~�c���x>�pЩ�U%`�l��w��@1�pTl�ro����x9�Yݢ�y�|�S�y�w\)�੍�sμ1N�#��-�L+M���i�6�2�%��@4mTR�D�M[R2'��y���#��ɢ�w�|Ou\[����߽!���H.�ذ(+᩼�_q����s\B|})�9�X��u���e�EA��(��_�~��+���fE�F�枽%��u�`�;���Z7~���1�P�/�	��#�(
��@��:�� �l?<]��{i��'\UE ���R�B��,��}0x�V��+6�w��Ur��̎j�3s����6{�K����Ӻ���Hd��x�������j�qA�d�ۛ���+U��Zi*O��h�F�i�$v5�)��h�?5(`P���.�S/�1��Fzp "��]����g� Ye�k�O3~d����{:�;1d市��
��6��É��M;�π���Hց�Z�a�Uؠ-0��Ky�ؖ�x9X���eK_Jl�G�@�
wD�X�E��Lf��K0@�VQ�G^�(�9:q���Q�i獈>Y`�s�Y� G|�D���|����F�h�2@A}R�')��*��4�����G4��4Sجޤ8�_�"��V����v+X�@��&�2}Gl��w�X���C�{+����u�8C��m�f���.d۬�&cZ�q!��b;S/����7ሸs��l�*L����Y���t���ʡÏ��݂&���YCX^��,��.̄�|���v�,7�bm��a#)���8��RC�*D���$�� �!D;�7���K�9'�PC��/��q�78��~���M/U��������z��W��Bvߡ��ш�=�Rq��0��6�@�Ɵ��.#���.M�@F�$��N��-����F �׬̖�jQQ���XaR��V[�ph�u��w�"$��&ǶS۶*��0B�ĵ?��*�y��� ��2�m���c�Ѕ���
b�Kﵬ������',�h_��Ȥ�W��Z���kI�i�MI��9}��RE�k�\
���v.��R�+u(��ߌL�����G�]�!,�e�.�y!s�+�U�/u������B�wc�����T�M�3D�A�/#��������bZ���Ǵ7�;6'�� nŢ~��m�j��|�U_� v�� _�x.8�DÙ��ʳ~=n.J��:�^�D�O/�͔���6��Sqr�����:|pX�����]���_��i& 3j�
�4���I�.�,5r#ʙaU]��'�d':���*���4�/k�m�O�G"r"��������s�bMD��J�Oa	c{I��L �vo*s��2��8$1V%��h����jT1�
�cv��qd-���nD1�+9�b��X��]v�Ω}�\+}�g���m<���r��_g��V�E����f���3�5�A+�P���7 {�t���.�K��V��i)0�t| �;c��e�Nn�fj!	U��z�ͭ �bWa\Q�s�P�k��� {�C����G��9����C~�c<��J4`��a��V��-d51��ɗ���ڎ��%�J�H�o��p��t�2�{���j.)�<�3{��d�^�T�7�3�*�G�UV�iwm�ؤP��E*i��뷞 s-���A?꾒�?%c��6�3��D���Q�3�d�A�H��5d#�I-P� �Gy<	$�Aj,LO{��S�Xs�?��*�/�k&����N�2$O�7���̶���6U���:�߶���>c��h���(����aǉ&j'n���H����/�%Qf"@�5s�ќQ��g=��S���|���|��U�����C�F�Q��l��LF�	��O u�+����2�w���0�x�4�S���1���?�1��J`�j��mT]q�f�nI}+�,���_��B3����pç?�~���CO�	��r�?>/z-��!غ�
��gW(�@�.� F���g�����?zKO���/8�[�Y��CZ�7����V��pb��}�S��^��D1��u�g��#��c�u���a�β"�:Q�e�T�!�ڢ�����i���,W12���'}։w����*��%i�uy��9Dج��{q1���+k{$���$ii�,D�d�J����:Py�%yd/�j�,��r�w��)��ҭ�Gn$f6�z�*�X�%�"xd���Y�P��Oϭ�XteW�~�.�9�(*�����Ⱦ�3{��Y�PY����`�81c�Cs{����uQ��4�
7U|md��ѫ���oSe��ϑB�@'?��
�.j���p��9D�^�Ӡ�˧�a�o�l%V�9�_�5f��a?|�%��]����ǐ`*��F�!��?�KZ��F�6
��`�:�Ű�[��]@�=؉�^���n���Yw�sH���g��� O�q�r	|!W���v���Tn��t�Yċe��e�	d;�Y���=�kO���!ν��R��b�t�5"�q��P�yzc3�@X�0��2�A� ��JWN��B�]�����+[�>t��Rr���lX>!��L���[�lU�á��@9]�H�͏;�$����p��Dit~�-+��):Q�����n���g�/��[^���6h������Χ��;'�m/S���_�zƓ,0�J�����Z��W�ϱ 3���8�,������<hplA�N	}����K��~�q�r���)́gFD��Y����ʧ��&�2C��

{%u��f���}j�]�x���-}9\��,�9HX6)��(�j�ׅV��q��V���`ME�^JP֎$�|��qD��#'� 5����Jz����sX��԰���*��&VAɀ����������%���"e|�5P�Ny�[��N��u쾱� �c�B��7v\���Q�ӌ�
���W[Y\�,��z����^��T0<u#.c͚��b�X�0�ixHa��4'���D���ʪ�騀a.UV��EI�e�#��tY��u�Bn/�u�[q���J������|��sԕ�/Q7�k���1*[�DG�s�&	4i����ߣ�I%�A0�,��S��;����g�u����첻EN_��A`�!��w�S,���(�)T-������m[�+@��b�@:t91�\��	c�8�Vk�>��(H��h�%�ے��eA�ک�-��2��##ހ�)},��`��ԋ�\�f>e �L�W8As��q?���LX2�y�w�7�hey M<yo$'h�݌��I�U��Y�ҭ�ɴ_�-��-I�n�����e0)�G�0}��M~���a�:k�y��g�k(�Q�%�Ќ)T�.���$uҬ_i�j8���g܎
���Y�Qd�z	���y@��<�E��Kډ�[.����\~���M�]�=!�4BZH�l������M�G�Ut��B�nV�j��YZX���w!b�cSt��噛�K�^��G	��p�H!fV�aG��w������&N(��5ߋ���<b�%�3�*�+�8�"iCV�4��l��7X�^rD3�UH�H7>��G�N�_DB_��?�E
L\�f>zI�>.�CD-�̐�-� XW�������;�����u��=��p��_k%8tV�0~����|��x�9h�im�������%$�HO;A�+yt$Ԍ�����t�� !wN����u@�e%
WO�� m4ǰ�fG��0}5/����X��tb��ޚ/;�Ov���{iӭ<�NOi��Q��űzE�t���$
�t��w��&:��-5��wl���F�y�#��CJ�rU��oҞ��c�}/ �h�����/<%W���aR�bq�NI�m�f���zm�*�~]XL\�x�=�<y���aK���D�9����W�\��?V�X���A�$S��^U�j;/������w#D�i�<J��|uޣ�Ta�k�c\�aR����^��*eH�uM�B����P�]3˘Ǽ Lx0���W�Y�(�c�'�Rgb�� ��yu]?�݆i9%؃�L��'b`�߀qhn3n�c`�N��������"�1Fm�.���a�u�V�Fc���� ���XlxV64EB    4b2f     d00�	`9'�%L���v����}�#���d�(7�Q��Y"܊�z���  oJ-",hP���M�*��U���Y��y����tY^W�Z��WF�.7��-�][��f��Db��5e=�IE�s�����I]	��M��w&5��9r��*��.���@R����(�_���0�]Q�wA��(]�����/���M��J6������CA�7�E0�� )�2ŚRY3��A���:�T�r�(UA��T���S�ǿ�VI-��'�o��74K^�%OF�y�Y�4�3�N�V� �|T�:���%L��=hޠ�}v.�X4����\Q�J�{�%(�Bi���"
���;�;�3��(���X��?�l8;�ۘ�#�`6�HL�o{����~r��Q"���Z�(����+��� +\��6�(�\"�-M��!�ҝ���ˑUjI����q	�����M$s�1�^g(�,7����t�d�hTU�_��	0�[&�@�w��=���n,6K&@�
7.~A���"d����?��(�4�(���uq��� ��r-I� o�qU�_��0u�[^��^a*}zσ� �p���e��n�����lN߬��?X2�N������1�~32�Ҝe����KE�S乣���|����}�@�P���P��O��j F�ge�	���h��Z���]:~���D���Q�h9���[F�6.��Wв��KO`}���,8���� :͕z���`)��v鄛Ƕm��6����x!g EPZ	k�M�+<�T�����/T������p+��_���e1��d�e��`ya�8��*Nm��u�ƍ$<�Ф��<�Y�詗�)��9�/�������u��{�(�ֺ5���NP�xb��R��7��S�T�Ci�q���d��(��Kh��&��=�~5��3(,I�^ �m7�
f���3-�A&+�y����>`i7a�2cd"7{m�a�1����0X<�2�B6{�I��/_Ye9�03l��jz����OH�U.�FR�"��kX�x">3�gj��!%\z:	m��6�̙�(�Y�I~��x���q����e���}�q/���͢"E�@U m|�lڿ��O����ٱ>�N�K1�6pK6��ds�K�&kKL��VT%S�� h���^*TK|jsCQ��̅��D��d�C�N�:7���댑G�sw9%���s�\������i\�N�LR�F�o7c�Z �VY�!�*��h��ڙ�ИoT�[�{!���U���^3|�pj^���;<��E_wr G3�i9��2��0�F{Md����#p�l�M����^.���S_+Jű�'��R�̍�'(C��vFM�r�d� ���g"��҃
7�++����	�����U��e;!�e ����g@f m���>eˬs���a("[v�4�%���i4��y�q߿���?*�HI?�/�47sC�rs-�x���������H�DJvms��~	L>XŜW�o�.WoNU���@�S�;ھyDp�(�9���}<]w.tZ�v16�I�O%)L�cg����{�çž�����?��mFy��6~s��>9��
�B��w�p��i0��4���1�w4�ĸ��~�Y�Μ�X�r
�å�l2�}�yJ��)�)8f�I{OS"A,�2p�>?�x/���tw�\5�����LCA�2��@��X�q�3xg.z-&ZdW�<$"H�f� ���Vft܈{�y?c��h�$��#�p �G3��E����IM�o+����L;��<�Ҝ`�ne�6��JVZv�tc+�F�&ly����?d�v�a�M���1>��mz��if�j���@��o�ެ����)Kyb����z8�)Q�%U���>�8�L��ݝNop��� �b�0�{dASJ��	������@<�"�;$��r�4�db�5-~o�6|�$��!����^,ˆ����X�S��,l�
Y�݆�SB���5)Rj���. ~�c�q\y�=՛��ß�x�����4QIgl]J߼��Ġ��g���:hW�O#�,Au�џn��uIj�W��e�q�,h���MD���Y�㗰}$P���73# �i����;U!F@�w��M<��ţ�۸�Fឱ�����Bq�Lf۰���N/~���&�.p�r}�N���RtWo%fײ��8$��պ-�&>'�>����
V���2Ӫ]nѷ��a�������=��чI6��7߮
�M�3��s���v�
5���%�������,d�u���Q|�-�}u����߰*2�Od�"�~�_QPQ���7�g@Np����uӟ�y\����P\C�I���
�GIt�Q���k$�[o% 6���$�f�~J�^�k9ߕ��{��c��y6��z��%�V#��G��R.��H] ��~�]�����.�֡3�tX�<�;w�̥��*��l)�T۝Ó�|��ШG�N�I ,��:�{�Q}����Q�>�!V4rX�:�Z�l��4�����jV`n�.ck).őI���v��f�,^2������sc�F�b*�5��݅�a!���<|mF�^�0��I[�fg�6��*p�o]#�|B���#�j5n!گ��q*O�`#g��e3/3�k��{OY����w����z���/"xo�[P+�Ũ6�p��'˖�A���oe�_��Hۛ*}�?�p3}I8a�1�7��.V��O�(AuCA�"�y0;�.�0<�<�,P��川�3������OF
C�Ow�/������|����Y�C8��o�I�q�f8�yN�M𘦃�o�.���	u��1�Cy�5���?����%=i�]��,CB$�̓IL�7D�:Xq'�m�=�s�G�j_��K�Ӫ0���A4�ԟ��qƇ[��@�u�7�/<I����+Rk������`������hEv�"�Y;K��-�Ն��^mJ[��R��	hGn?�ȩ� PҔ���{`�lD�=<�pΣ�
yh��&BRxD���y����;%��p|ycL�����f} u�;�0��7~4�[��..����$�� 6"��:F�Pe�N_���x:�9|}���za:3NkV���y�*�pV(��U��s�&.��K�ݬY�+��.ڢ����BQ��|�����MO�E�3�H	ª �f۵��x|���$Zy.�e7UI��ڔ~-_+�=�+���nH�.����	�Sv���K�*]��B$��"���P��IH�i�{���Z=W