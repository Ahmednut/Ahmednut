XlxV64EB    24ab     c50UJ�?_��X�Գg&J<�9+�M��v�ȱ��o���f?��D]n��r�<���[@�	oE�(b�[�]E���\���N�}��6�N%P��L�mlL�s6v7[�[>L�b%B�ݝ��ż�f����q��E�C��I��o���n�`��<^c>d�W�??&���Ni)d)���ͮ	��YO̶��m:%�00�j3!��F��߱7m�X�	k˺w[ B)!/�JAE�J�z�M	5�/6d�M3䡾���$��(pmF╸+������[��XyOM���Ii�cϡS`9�$^A�ȅ9���;�)�^w�W����VH_�}U��#�)o���]�b����%��#�$�Z]y�욫�RxV}7L"' \%��{Tm�����Hh�kCM_,�&Ksm<yI���<���S�\B�)6�W�`݋���W��a��EM�ɗ�Lˍ��W+�1v���g��c�EB:�~�DD�����P�����u�K�^�I�:�L��@1�p�!��(3>/Et���&n��U�83tͪ���bm��XrDG3���݋^\����C�b!�*f��mM���ae�J}=���Q��/H4ӓ���\�}��{�?��:�S[BB}l%S�~. �>P�%�q;jV}��x�(p͖����gby�R��?Xj������UĻnGd��%kvm�c�@<Q�h��cﻺi�p�Q��ZCanv�Ջ�`B?[�*/�����t�-1�R���e|�Փ_�t{2*��=�]k�&�m-��C�J�a܏�$��{6��E�N=��$oQT;N�R)��l3#ҏ��tJ;7�t�R@�P`�c���IA����{�_��/���[:e�M�2�M��� �ꄶ�w�=�{�	�"�FP4'�F��I��R���Wu�(�{�� ƨ�w6'�7I,��=��E\��5������*�{p^|�-�P��fˢ�"�G}#���}�GL�ꝸ0p������2�+���#�U�s����F�t[�M4�(װ0��7ۆlu��E�ФС��`�\�}g�n��
�N��\�پm���k�*���X|�����[�J����?�ZgPa%�_�n˝u}�WyֽЅ�<ԵK� ��#�<�8�X�Y�΂SS�f�@�Hh<�$;�0�zt[��F9_W��W�*�7�h����!B�(#RS�WF��r�b��*9�_�"�=�m���m̚uh������Z�9��c:N��B���-t���=��GE�~8r�5gAD:�a��x��S~�;�YR�I�`��E��ݟ�Ñc|�ٟT5���X�&�$��=�{��z1�
SS�l%��2���M��H�š����Q�*�N����c���q�k�������Y��4˧\� �u`�?e�5`_�����k��_G�*"<�X��
o\���nMyIK�su�
y��U���÷w���g��\�k=5�E71=�L/�Hb�������
����L'N�Ѽ���γ�/>�I�T��"F6��%��@[�Rm���:^ˎ�풟�OĐ��L����q�S�Zy�]�s�A��(������l��܊B��]���jآ.��`ƲD�/)f�<׹LR���i$�`qL���rSнfP�#�<��:���n�"S���'��ie�?�R�sFuS_������W����,^
A������\����"]��mB�Z��
��;��!�M���:��<�����S�����f��z��ހݧ�y�@]Í��m��ЗH�v�Q��N"��U*$���\�0"c#�#Z�;���%gb`L�x�x)<`�����R�*��%r[��	�ͺ����RM*h'����}�ȹ[&lOv�G���е��f�[.@������4
f]�h@��T k^[���Q���,�EY4ƪ�wW���2��79�P�:x_��I��̱��4nnRn�b����|�K(�+�`����*W�t�h>�Yx�@�1��W��: !'dЖPICbKb?� S��
]��㷥��GLI��?�KLʁm{[K���F���?�_�������;���\��H�S�):�T�do��&��%9ʰMDi9�)��� ��p�IWl؆�5�"	|r�Xھ�c��휘F-�L��$��׶�14��C���5:,����O�[M]rߡS��s���v��c��<Ǵ7[�c�w.S7�
���1�S������eU��gM|8!��0���!��Ŧ=�}������*I�HɣӋ|�%��c�-��:阘4��3b�"�,�.Z���];����v�S�H2�X5��l�N7�#�pB(ɵ����Ĳ�R�؞�2�ݳ9>�ə�5���Q��F�'evS՝Q�	n��e�QH��Aq^ڊ��M����s�緋�B���ݓ��,+SI��-�} �͌�|G�Ղ��>�M��m�66�۠�͟��P�0(�bY)2�w'���U��nr�߿z3{��c=�ރk�ZvNAݠJ�z�� A�o2zK��S�e�Au��@J����g�|M:�ma#�0֐-�������z�)S�4��\ �����~jV��M
�aCu���2u�
�#�29�k�~Q���y+�sU��3�;�.R���:E���م; A���?�<;oV�����@�����vY<<��9��TQp���5w�f���?�٫@&���x�(���_��-n��.evFx,�6�������nH}�tڴr���>T�o��� H�5gVzw. x�u���}|������]R=\�����S�J���с�[��~�d�5�ktL���O����w����u�Q���M+L�1xAT���,m�P<@�e�hWV�vh�����P�[����V^�1��mГ�01��|���a�tV!ؠB�[�1��GyB�X]�Ȇ�G���3�D�r�r��*oMş,é������ݼ�͑��rt
_T7o�L��-a�_,�m�C��>N~-��q�Li���	�S] R����t�&��R*a�K`k���Q��k:;���[l�.t�,�,�7�iِF��"�"�����s lЯ��h��������m�6::��,��Q����Zq�}��