--------------------------------------------------------------------------------
--
--    ****                              *
--   ******                            ***
--   *******                           ****
--   ********    ****  ****     **** *********    ******* ****    ***********
--   *********   ****  ****     **** *********  **************  *************
--   **** *****  ****  ****     ****   ****    *****    ****** *****     ****
--   ****  ***** ****  ****     ****   ****   *****      ****  ****      ****
--  ****    *********  ****     ****   ****   ****       ****  ****      ****
--  ****     ********  ****    *****  ****    *****     *****  ****      ****
--  ****      ******   ***** ******   *****    ****** *******  ****** *******
--  ****        ****   ************    ******   *************   *************
--  ****         ***     ****  ****     ****      *****  ****     *****  ****
--                                                                       ****
--          I N N O V A T I O N  T O D A Y  F O R  T O M M O R O W       ****
--                                                                        ***
--
--------------------------------------------------------------------------------
-- File        : $Id: lyt_idelayctrl.vhd,v 1.1 2015/04/10 19:48:37 sqa Exp $
--------------------------------------------------------------------------------
-- Description :
--------------------------------------------------------------------------------
-- Notes / Assumptions :
--------------------------------------------------------------------------------
-- Copyright (c) 2012 Nutaq inc.
--------------------------------------------------------------------------------
-- $Log: lyt_idelayctrl.vhd,v $
-- Revision 1.1  2015/04/10 19:48:37  sqa
-- bas first commit
--
-- Revision 1.1  2013/10/22 13:30:25  julien.roy
-- Add idelayctrl core
--
--
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library unisim;
  use unisim.vcomponents.all;

entity lyt_idelayctrl is
    port
    (
        i_rst_p       : in  std_logic;
        i_clk_p       : in  std_logic;
        o_rdy_p       : out std_logic
    );
end entity lyt_idelayctrl;

------------------------------------------------------------------------------
-- Architecture section
------------------------------------------------------------------------------
architecture arch of lyt_idelayctrl is

begin

  -- IDELAYCTRL instance
  idelayctrl_inst : IDELAYCTRL
    port map (
      RDY 	 => o_rdy_p,
      REFCLK => i_clk_p,
      RST 	 => i_rst_p
    );

end arch;
