XlxV64EB    1fe1     ad0�����7&���#{��ӱW7R��b�h�6~b�m�t�5�::���B�a�2�$�������X�a(n�̊��U$g�#����#��:朲(	Aҥ.�η���EvH�ܤq� -���ǯ$]�	)��l�YѐԲ�k�E�,<���}Ŝ��S�x,C� �������%�q��׬D�I�q�Ak�fH�Sj��\m�	����ar1�� dQD�Ք�	1�~U��ehw��h�����
V(ՕAޓ�Qmv�,�, �p��X9q�b�_ � �.�LQ_���t%	B��3�1S�VzN��Pk�է��O'0fe�%L$�L\9㛖��u�Gq R�+�����s���]:��1'�{��WF�{��̸�ܔ'(^f�t� �-z�C���I�^s�$�!|z?��"MF��#�c���!2�g�<��啓��+����
��H�L
,����S�4鱎{�
z��H%�Pr�e��O>J��*�n�b��&��;΍�J��z˒��e_S^r�4l;.ྡM\�v���D:�󓂸��0��nq<���h�\]�9`П8�k�k[X%1Oڂ@	�� �b�ET�|\#&m�r�>`��[�
�Zf�����E#�/�^���N�������}�8��C�5��u����yyX=��0��j�i��� �t�>
���k�G��A�38H�l��O3g#���$��S�V{�LvBD�L��g���۪o�@w�U>9�嗀`�&^N�:0"�|����)��ĭ���aE���[�H+�)�$�Ù���N�*���+eX��,)�l���Mu��L$��k l 
�|��_���D�_;�b��Td������b �2�按$&�\��,���`�o	?�;�+�6��}C�T� �b�,���1��/��[��i�C@hJq���ծ#ϗ�MCԊ���؜b����iN��Լo���T̞}/���c�@��Ft.0ґ.��,����*�`h�cVB�Em{V1���,���ɸ�{�U��;~uc�Q��*c�a���t��P|t�&!�t�%�\4j4;G����o�*�<��6��ْ��&�4���|�/v�s�r��.~: ɛ��2�D��jz���& ���y�gR^Q�Ks=��;���#1̟rnAAKmW���I�$�{B��Ž��^�>YR����ʔ"@h�)�l7�
� ���j,�Vk��c}�یQ�2�'ο,�TyJ���тr��H�^ A7�@%����`��'���s��N1��|i��ǟ�^>=R+ٍMB�#�'�3�:�%Ԯ^�+7L�h6�c!u'�iJe������>���E0�~fZҖ��������4j���8�Z��%�W�H����������������J��2ϡ��'6��˃@���(��OLn�6�V�@��V��U��r5Ĭ�	����?�d6�>#�[�V�~�,�
W!�+sD�l���E�\s�3`��мi0�r��$�J�L��c_�-�����ؓW�
��rq�F�t!ԃ��̆�z&��S�������
�4��b������/��Xq�	�{|΋Q�G&���ڑN.$�����`ۅ��2�¸<9 ���\x�J㥏t\ۮcJ�"8�l�Z�(�p4��*M�]���{䜱�w��z*��A����A��d��H/�`�!@ӝwTF(P��0`�|S���	u1���f�_�>Ӹ�i�϶\�������uyx5&��p���B��{Q�bY6S���	��c"?�x���)���#���Ѻ�ogL�_�5��� �-C��v�C��ϩ-��<�����5!gJ�A=���tl����r�L�ju>��:�_"�����C�!�S@��X�3�33E�$�y�������o�dV��I��B
R�%�cqd�Rtqu�QI����V�=�� \�h��R�p�篹���"I�J�.���Q%�����<���	�C@Qsƚp3�Q:���o������������I��,vT��XhǺ���L��`�i"��i�EX��v���A7�U��Q!���i����^��4S���R��}P74̩i��=�i���f�~}�:=#��re4+m�=�!֩�Je�ù"lq�+�$(F^�������R!-?�;�!h:2�6�K	�^��|̲Ȣ����{y>>���r��Q`�d�u��Hn�J�K�^�ci�P�n�}G-�?�Mn)P-���q�%_ކN^�(T"��%��FǬ�Y�cAKÍ�ZH�0<��8����Q/���n.s����d��x���7'|�>�#V?˾��>46|
��M<�Tɧ��'�U��ò%:�+I�2��Q�vVIt�k��]�GK��bT�R�+�NO��5�r>v�
}3�Z��_�2c�?b���e<_�d���-e�%m�f��o�-�V��������VѮd�MrX(�pVΛ�ő��_Z��U.��=2ڕ+@�[�+�D�K"��p/p��Z%�Ni���K3�+a|����D�#�5U�k�6Et�d�t�ڣ`�Ė��'�0�-F���uAi��cf�0)Ҵ����b��f��t/���w��{���m�������8u6��R}n~��}3���P��7�����f��Ř��'7R ckh�Jm���_U>�Xu�`O�M��J�XO֑'[�do%���Ź�̮s/���%گ��,B)ї�= a�!)&�,�z_���[��2{�