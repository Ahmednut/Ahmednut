--------------------------------------------------------------------------------
--
--    ****                              *
--   ******                            ***
--   *******                           ****
--   ********    ****  ****     **** *********    ******* ****    ***********
--   *********   ****  ****     **** *********  **************  *************
--   **** *****  ****  ****     ****   ****    *****    ****** *****     ****
--   ****  ***** ****  ****     ****   ****   *****      ****  ****      ****
--  ****    *********  ****     ****   ****   ****       ****  ****      ****
--  ****     ********  ****    *****  ****    *****     *****  ****      ****
--  ****      ******   ***** ******   *****    ****** *******  ****** *******
--  ****        ****   ************    ******   *************   *************
--  ****         ***     ****  ****     ****      *****  ****     *****  ****
--                                                                       ****
--          I N N O V A T I O N  T O D A Y  F O R  T O M M O R O W       ****
--                                                                        ***
--
--------------------------------------------------------------------------------
-- Filename:          user_logic.vhd
-- Version:           v1_00_a
-- Description:       User Logic implementation module
-- Generated by:      julien.roy
-- Date:              2013-01-04 13:33:18
-- Generated:         using LyrtechRD REGGENUTIL based on Xilinx IPIF Wizard.
-- VHDL Standard:     VHDL'93
------------------------------------------------------------------------------
-- Copyright (c) 2001-2012 LYRtech RD Inc.  All rights reserved.
------------------------------------------------------------------------------
--
-----------------------------------------------------------------------------
-- Register Memory Map & Description
-----------------------------------------------------------------------------
-- BASEADDR + 0x0   INFO    ADAC250 Core ID and Version
--   15:0 Version R
--   31:16 CoreID R

-- BASEADDR + 0x4   ADCCTRL    Drive ADC's based signal
--   14:10 TriggerDelay R W O=ov5_TriggerDelay_p
--   15:15 CoreResetPulse P O=o_CoreResetPulse_p
--   1:0 AdcRun R W O=ov2_AdcRun_p
--   31:16 rsvd2 R
--   3:2 AdcStart R W O=ov2_AdcStart_p
--   4:4 AdcDataFormat R W O=o_AdcDataFormat_p
--   5:5 AdcSpiReset R W O=o_AdcSpiReset_p
--   6:6 ADCAOvr R I=i_ADCAOvr_p
--   7:7 rsvd1 R
--   8:8 ADCBOvr R I=i_ADCBOvr_p
--   9:9 AdcResetMmcm R W O=o_AdcResetMmcm_p

-- BASEADDR + 0x8   DACCTRL    Drive DAC's based signal
--   0:0 DacReset R W O=o_DacReset_p
--   1:1 DacDataClkLocked R I=i_DacDataClkLocked_p
--   31:8 rsvd2 R
--   4:2 DacAMuxSelect R W O=ov3_DacAMuxSelect_p
--   7:5 DacBMuxSelect R W O=ov3_DacBMuxSelect_p

-- BASEADDR + 0xc   MISCCTRL    Drive clock pll 's based signal
--   0:0 PllStatus R I=i_PllStatus_p
--   1:1 PllFunction R W O=o_PllFunction_p
--   10:10 UpdaterBusy R I=i_UpdaterBusy_p
--   11:11 SpiBusy R I=i_SpiBusy_p
--   12:12 SpiReq R W O=o_SpiReq_p
--   13:13 SpiGnt R I=i_SpiGnt_p
--   14:14 SpiAck R I=i_SpiAck_p
--   2:2 ClkMuxConfig R W O=o_ClkMuxConfig_p
--   3:3 ClkMuxLoad R W O=o_ClkMuxLoad_p
--   31:15 rsvd R
--   5:4 ClkMuxSin R W O=ov2_ClkMuxSin_p
--   7:6 ClkMuxSout R W O=ov2_ClkMuxSout_p
--   9:8 RSVD1 R W

-- BASEADDR + 0x10   SPI0    Spi reg 0

-- BASEADDR + 0x14   SPI1    Spi reg 1

-- BASEADDR + 0x18   SPI2    Spi reg 2

-- BASEADDR + 0x1c   SPI3    Spi reg 3

-- BASEADDR + 0x20   SPI4    Spi reg 4

-- BASEADDR + 0x24   SPI5    Spi reg 5

-- BASEADDR + 0x28   SPI6    Spi reg 6

-- BASEADDR + 0x2c   SPI7    Spi reg 7

-- BASEADDR + 0x30   SPI8    Spi reg 8

-- BASEADDR + 0x34   ADCDELAYCTRL    Control ADC data and clock input delays
--   10:10 AdcPatternError R I=i_AdcPatternError_p
--   31:11 rsvd R
--   4:0 AdcIdelayValue R W O=ov5_AdcIdelayValue_p
--   9:5 AdcClkIdelayValue R W O=ov5_AdcClkIdelayValue_p

-- BASEADDR + 0x38   DACDELAYCTRL    Control DAC data and clock output delays
--   31:10 rsvd R
--   4:0 DacIdelayValue R W O=ov5_DacIdelayValue_p
--   9:5 DacClkIdelayValue R W O=ov5_DacClkIdelayValue_p

-- BASEADDR + 0x3c   FREQCNTCLK    Clock frequency counter control and status
--   15:0 FreqCntClkCnt R I=iv16_FreqCntClkCnt_p
--   17:16 FreqCntClkSel R W O=ov2_FreqCntClkSel_p
--   31:18 rsvd R

--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library proc_common_v3_00_a;
use proc_common_v3_00_a.proc_common_pkg.all;

-- DO NOT EDIT ABOVE THIS LINE --------------------

--USER libraries added here

------------------------------------------------------------------------------
-- Entity section
------------------------------------------------------------------------------
-- Definition of Generics:
--   C_NUM_REG                    -- Number of software accessible registers
--   C_SLV_DWIDTH                 -- Slave interface data bus width
--
-- Definition of Ports:
--   Bus2IP_Clk                   -- Bus to IP clock
--   Bus2IP_Resetn                -- Bus to IP reset
--   Bus2IP_Data                  -- Bus to IP data bus
--   Bus2IP_BE                    -- Bus to IP byte enables
--   Bus2IP_RdCE                  -- Bus to IP read chip enable
--   Bus2IP_WrCE                  -- Bus to IP write chip enable
--   IP2Bus_Data                  -- IP to Bus data bus
--   IP2Bus_RdAck                 -- IP to Bus read transfer acknowledgement
--   IP2Bus_WrAck                 -- IP to Bus write transfer acknowledgement
--   IP2Bus_Error                 -- IP to Bus error response
------------------------------------------------------------------------------

entity user_logic is
  generic
  (
    -- ADD USER GENERICS BELOW THIS LINE ---------------
    --USER generics added here
    -- ADD USER GENERICS ABOVE THIS LINE ---------------

    -- DO NOT EDIT BELOW THIS LINE ---------------------
    -- Bus protocol parameters, do not add to or delete
    C_NUM_REG                      : integer              := 16;
    C_SLV_DWIDTH                   : integer              := 32
    -- DO NOT EDIT ABOVE THIS LINE ---------------------
  );
  port
  (
    -- ADD USER PORTS BELOW THIS LINE ------------------
    --USER ports added here
    -- ADD USER PORTS ABOVE THIS LINE ------------------
    -- User ports
    i_CoreReset_p : in std_logic;

    ov5_TriggerDelay_p : out std_logic_vector(4 downto 0);
    o_CoreResetPulse_p : out std_logic;
    ov2_AdcRun_p : out std_logic_vector(1 downto 0);
    ov2_AdcStart_p : out std_logic_vector(1 downto 0);
    o_AdcDataFormat_p : out std_logic;
    o_AdcSpiReset_p : out std_logic;
    i_ADCAOvr_p : in std_logic;
    i_ADCBOvr_p : in std_logic;
    o_AdcResetMmcm_p : out std_logic;
    o_DacReset_p : out std_logic;
    i_DacDataClkLocked_p : in std_logic;
    ov3_DacAMuxSelect_p : out std_logic_vector(2 downto 0);
    ov3_DacBMuxSelect_p : out std_logic_vector(2 downto 0);
    i_PllStatus_p : in std_logic;
    o_PllFunction_p : out std_logic;
    i_UpdaterBusy_p : in std_logic;
    i_SpiBusy_p : in std_logic;
    o_SpiReq_p : out std_logic;
    i_SpiGnt_p : in std_logic;
    i_SpiAck_p : in std_logic;
    o_ClkMuxConfig_p : out std_logic;
    o_ClkMuxLoad_p : out std_logic;
    ov2_ClkMuxSin_p : out std_logic_vector(1 downto 0);
    ov2_ClkMuxSout_p : out std_logic_vector(1 downto 0);
    ov9_SpiWriteaddr_p : out std_logic_vector(8 downto 0);
    ov9_SpiReadaddr_p : out std_logic_vector(8 downto 0);
    ov32_SpiDin_p : out std_logic_vector(31 downto 0);
    iv32_SpiDout_p : in std_logic_vector(31 downto 0);
    i_AdcPatternError_p : in std_logic;
    ov5_AdcIdelayValue_p : out std_logic_vector(4 downto 0);
    ov5_AdcClkIdelayValue_p : out std_logic_vector(4 downto 0);
    ov5_DacIdelayValue_p : out std_logic_vector(4 downto 0);
    ov5_DacClkIdelayValue_p : out std_logic_vector(4 downto 0);
    iv16_FreqCntClkCnt_p : in std_logic_vector(15 downto 0);
    ov2_FreqCntClkSel_p : out std_logic_vector(1 downto 0);
    -- Bus protocol ports, do not add to or delete
    Bus2IP_Clk                     : in  std_logic;
    Bus2IP_Resetn                  : in  std_logic;
    Bus2IP_Data                    : in  std_logic_vector(C_SLV_DWIDTH-1 downto 0);
    Bus2IP_BE                      : in  std_logic_vector(C_SLV_DWIDTH/8-1 downto 0);
    Bus2IP_RdCE                    : in  std_logic_vector(C_NUM_REG-1 downto 0);
    Bus2IP_WrCE                    : in  std_logic_vector(C_NUM_REG-1 downto 0);
    IP2Bus_Data                    : out std_logic_vector(C_SLV_DWIDTH-1 downto 0);
    IP2Bus_RdAck                   : out std_logic;
    IP2Bus_WrAck                   : out std_logic;
    IP2Bus_Error                   : out std_logic
  );

 attribute MAX_FANOUT : string;
 attribute SIGIS : string;
 attribute SIGIS of Bus2IP_Clk    : signal is "CLK";
 attribute SIGIS of Bus2IP_Resetn : signal is "RST";

end entity user_logic;

------------------------------------------------------------------------------
-- Architecture section
------------------------------------------------------------------------------

architecture IMP of user_logic is

-------------------------------------------------------------------------------
-- Constant declarations
-------------------------------------------------------------------------------


-------------------------------------------------------------------------------
--     ************** Function declaratin *******************                   
-- Return a std_logic_vector with only one bit set to one.
-- The argument BitPosition represent the bit position to set to one, starting with 0.
-- The argument Width represent the width of the returned std_logic_vector.
-------------------------------------------------------------------------------
  function OneHotVector( BitPosition : integer;                              
                Width : integer)                                             
                return std_logic_vector                                      
  is                                                                         
    variable Result                   : std_logic_vector(Width - 1 downto 0);

  begin                        
    Result := (others => '0'); 
    Result(BitPosition) := '1';
    return Result;             
  end OneHotVector;            
-------------------------------------------------------------------------------
-- Signal and Type Declarations
-------------------------------------------------------------------------------

  signal v5_TriggerDelay_s                     : std_logic_vector(4 downto 0);
  signal CoreResetPulse_s                     : std_logic;
  signal v2_AdcRun_s                     : std_logic_vector(1 downto 0);
  signal v2_AdcStart_s                     : std_logic_vector(1 downto 0);
  signal AdcDataFormat_s                     : std_logic;
  signal AdcSpiReset_s                     : std_logic;
  signal AdcResetMmcm_s                     : std_logic;
  signal DacReset_s                     : std_logic;
  signal v3_DacAMuxSelect_s                     : std_logic_vector(2 downto 0);
  signal v3_DacBMuxSelect_s                     : std_logic_vector(2 downto 0);
  signal PllFunction_s                     : std_logic;
  signal SpiReq_s                     : std_logic;
  signal ClkMuxConfig_s                     : std_logic;
  signal ClkMuxLoad_s                     : std_logic;
  signal v2_ClkMuxSin_s                     : std_logic_vector(1 downto 0);
  signal v2_ClkMuxSout_s                     : std_logic_vector(1 downto 0);
  signal v2_RSVD1_s                     : std_logic_vector(1 downto 0);
  signal v5_AdcIdelayValue_s                     : std_logic_vector(4 downto 0);
  signal v5_AdcClkIdelayValue_s                     : std_logic_vector(4 downto 0);
  signal v5_DacIdelayValue_s                     : std_logic_vector(4 downto 0);
  signal v5_DacClkIdelayValue_s                     : std_logic_vector(4 downto 0);
  signal v2_FreqCntClkSel_s                     : std_logic_vector(1 downto 0);
  signal slv_reg_write_sel              : std_logic_vector(15 downto 0);
  signal slv_reg_read_sel               : std_logic_vector(15 downto 0);
  signal slv_ip2bus_data                : std_logic_vector(C_SLV_DWIDTH-1 downto 0);
  signal slv_read_ack                   : std_logic;
  signal slv_write_ack                  : std_logic;

------------------------------------------------------------------------------
begin
------------------------------------------------------------------------------

-------------------------------------------------------------------------------
-- Begin architecture
-------------------------------------------------------------------------------

-- swap bits
WrCeBitSwap: for i in 0 to slv_reg_write_sel'high generate
  slv_reg_write_sel(i) <= Bus2IP_WrCE(slv_reg_write_sel'high - i);
end generate WrCeBitSwap;

RdCeBitSwap: for i in 0 to slv_reg_read_sel'high generate
  slv_reg_read_sel(i)  <= Bus2IP_RdCE(slv_reg_read_sel'high - i);
end generate RdCeBitSwap;

-- generate write/read ack
  slv_write_ack <=   Bus2IP_WrCE(0) or   Bus2IP_WrCE(1) or   Bus2IP_WrCE(2) or   Bus2IP_WrCE(3) or   Bus2IP_WrCE(4) or   Bus2IP_WrCE(5) or   Bus2IP_WrCE(6) or   Bus2IP_WrCE(7) or   Bus2IP_WrCE(8) or   Bus2IP_WrCE(9) or   Bus2IP_WrCE(10) or   Bus2IP_WrCE(11) or   Bus2IP_WrCE(12) or   Bus2IP_WrCE(13) or   Bus2IP_WrCE(14) or   Bus2IP_WrCE(15);
  slv_read_ack  <=   Bus2IP_RdCE(0) or   Bus2IP_RdCE(1) or   Bus2IP_RdCE(2) or   Bus2IP_RdCE(3) or   Bus2IP_RdCE(4) or   Bus2IP_RdCE(5) or   Bus2IP_RdCE(6) or   Bus2IP_RdCE(7) or   Bus2IP_RdCE(8) or   Bus2IP_RdCE(9) or   Bus2IP_RdCE(10) or   Bus2IP_RdCE(11) or   Bus2IP_RdCE(12) or   Bus2IP_RdCE(13) or   Bus2IP_RdCE(14) or   Bus2IP_RdCE(15);

 -- implement slave model software accessible register(s)
 SLAVE_REG_WRITE_PROC : process( Bus2IP_Clk ) is
 begin

  if Bus2IP_Clk'event and Bus2IP_Clk = '1' then
    if Bus2IP_Resetn = '0' then
      v5_TriggerDelay_s <= "00000";
      CoreResetPulse_s <= '0';
      v2_AdcRun_s <= "00";
      v2_AdcStart_s <= "00";
      AdcDataFormat_s <= '0';
      AdcSpiReset_s <= '0';
      AdcResetMmcm_s <= '0';
      DacReset_s <= '0';
      v3_DacAMuxSelect_s <= "000";
      v3_DacBMuxSelect_s <= "000";
      PllFunction_s <= '0';
      SpiReq_s <= '0';
      ClkMuxConfig_s <= '0';
      ClkMuxLoad_s <= '0';
      v2_ClkMuxSin_s <= "00";
      v2_ClkMuxSout_s <= "00";
      v2_RSVD1_s <= "00";
      v5_AdcIdelayValue_s <= "10000";
      v5_AdcClkIdelayValue_s <= "00000";
      v5_DacIdelayValue_s <= "00000";
      v5_DacClkIdelayValue_s <= "00000";
      v2_FreqCntClkSel_s <= "00";

    else

  -- Synchronous reset
  if ( i_CoreReset_p = '1' ) then
    v5_TriggerDelay_s <= "00000";
    CoreResetPulse_s <= '0';
    v2_AdcRun_s <= "00";
    v2_AdcStart_s <= "00";
    AdcDataFormat_s <= '0';
    AdcSpiReset_s <= '0';
    AdcResetMmcm_s <= '0';
    DacReset_s <= '0';
    v3_DacAMuxSelect_s <= "000";
    v3_DacBMuxSelect_s <= "000";
    PllFunction_s <= '0';
    SpiReq_s <= '0';
    ClkMuxConfig_s <= '0';
    ClkMuxLoad_s <= '0';
    v2_ClkMuxSin_s <= "00";
    v2_ClkMuxSout_s <= "00";
    v2_RSVD1_s <= "00";
    v5_AdcIdelayValue_s <= "10000";
    v5_AdcClkIdelayValue_s <= "00000";
    v5_DacIdelayValue_s <= "00000";
    v5_DacClkIdelayValue_s <= "00000";
    v2_FreqCntClkSel_s <= "00";
  end if;

  CoreResetPulse_s <= '0';
      case slv_reg_write_sel is

        when OneHotVector(1,16) =>
          if (Bus2IP_BE(1) = '1') then
            v5_TriggerDelay_s <= Bus2IP_Data(14 downto 10);
          end if;
          if (Bus2IP_BE(1) = '1') then
            CoreResetPulse_s <= Bus2IP_Data(15);
          end if;
          if (Bus2IP_BE(0) = '1') then
            v2_AdcRun_s <= Bus2IP_Data(1 downto 0);
          end if;
          if (Bus2IP_BE(0) = '1') then
            v2_AdcStart_s <= Bus2IP_Data(3 downto 2);
          end if;
          if (Bus2IP_BE(0) = '1') then
            AdcDataFormat_s <= Bus2IP_Data(4);
          end if;
          if (Bus2IP_BE(0) = '1') then
            AdcSpiReset_s <= Bus2IP_Data(5);
          end if;
          if (Bus2IP_BE(1) = '1') then
            AdcResetMmcm_s <= Bus2IP_Data(9);
          end if;

        when OneHotVector(2,16) =>
          if (Bus2IP_BE(0) = '1') then
            DacReset_s <= Bus2IP_Data(0);
          end if;
          if (Bus2IP_BE(0) = '1') then
            v3_DacAMuxSelect_s <= Bus2IP_Data(4 downto 2);
          end if;
          if (Bus2IP_BE(0) = '1') then
            v3_DacBMuxSelect_s <= Bus2IP_Data(7 downto 5);
          end if;

        when OneHotVector(3,16) =>
          if (Bus2IP_BE(0) = '1') then
            PllFunction_s <= Bus2IP_Data(1);
          end if;
          if (Bus2IP_BE(1) = '1') then
            SpiReq_s <= Bus2IP_Data(12);
          end if;
          if (Bus2IP_BE(0) = '1') then
            ClkMuxConfig_s <= Bus2IP_Data(2);
          end if;
          if (Bus2IP_BE(0) = '1') then
            ClkMuxLoad_s <= Bus2IP_Data(3);
          end if;
          if (Bus2IP_BE(0) = '1') then
            v2_ClkMuxSin_s <= Bus2IP_Data(5 downto 4);
          end if;
          if (Bus2IP_BE(0) = '1') then
            v2_ClkMuxSout_s <= Bus2IP_Data(7 downto 6);
          end if;
          if (Bus2IP_BE(1) = '1') then
            v2_RSVD1_s <= Bus2IP_Data(9 downto 8);
          end if;

        when OneHotVector(13,16) =>
          if (Bus2IP_BE(0) = '1') then
            v5_AdcIdelayValue_s <= Bus2IP_Data(4 downto 0);
          end if;
          if (Bus2IP_BE(0) = '1') then
            v5_AdcClkIdelayValue_s(2 downto 0) <= Bus2IP_Data(7 downto 5);
          end if;
          if (Bus2IP_BE(1) = '1') then
            v5_AdcClkIdelayValue_s(4 downto 3) <= Bus2IP_Data(9 downto 8);
          end if;

        when OneHotVector(14,16) =>
          if (Bus2IP_BE(0) = '1') then
            v5_DacIdelayValue_s <= Bus2IP_Data(4 downto 0);
          end if;
          if (Bus2IP_BE(0) = '1') then
            v5_DacClkIdelayValue_s(2 downto 0) <= Bus2IP_Data(7 downto 5);
          end if;
          if (Bus2IP_BE(1) = '1') then
            v5_DacClkIdelayValue_s(4 downto 3) <= Bus2IP_Data(9 downto 8);
          end if;

        when OneHotVector(15,16) =>
          if (Bus2IP_BE(2) = '1') then
            v2_FreqCntClkSel_s <= Bus2IP_Data(17 downto 16);
          end if;
        when others =>
          null;
      end case;
    end if;
  end if;

 end process SLAVE_REG_WRITE_PROC;

 -- implement slave model software accessible register(s) read mux
SLAVE_REG_READ_PROC : process( iv32_SpiDout_p, v5_TriggerDelay_s, slv_reg_read_sel, v2_AdcRun_s, v2_AdcStart_s, AdcDataFormat_s, AdcSpiReset_s, i_ADCAOvr_p, i_ADCBOvr_p, AdcResetMmcm_s, DacReset_s, i_DacDataClkLocked_p, v3_DacAMuxSelect_s, v3_DacBMuxSelect_s, i_PllStatus_p, PllFunction_s, i_UpdaterBusy_p, i_SpiBusy_p, SpiReq_s, i_SpiGnt_p, i_SpiAck_p, ClkMuxConfig_s, ClkMuxLoad_s, v2_ClkMuxSin_s, v2_ClkMuxSout_s, v2_RSVD1_s, v5_AdcIdelayValue_s, v5_AdcClkIdelayValue_s, i_AdcPatternError_p, v5_DacIdelayValue_s, v5_DacClkIdelayValue_s, iv16_FreqCntClkCnt_p, v2_FreqCntClkSel_s) is
 begin
   case slv_reg_read_sel is

        when OneHotVector(0,16) =>
          slv_ip2bus_data(15 downto 0) <= X"0200";
          slv_ip2bus_data(31 downto 16) <= X"A250";

        when OneHotVector(1,16) =>
          slv_ip2bus_data(14 downto 10) <= v5_TriggerDelay_s;
          slv_ip2bus_data(1 downto 0) <= v2_AdcRun_s;
          slv_ip2bus_data(31 downto 16) <= "0000000000000000";
          slv_ip2bus_data(3 downto 2) <= v2_AdcStart_s;
          slv_ip2bus_data(4) <= AdcDataFormat_s;
          slv_ip2bus_data(5) <= AdcSpiReset_s;
          slv_ip2bus_data(6) <= i_ADCAOvr_p;
          slv_ip2bus_data(7) <= '0';
          slv_ip2bus_data(8) <= i_ADCBOvr_p;
          slv_ip2bus_data(9) <= AdcResetMmcm_s;

        when OneHotVector(2,16) =>
          slv_ip2bus_data(0) <= DacReset_s;
          slv_ip2bus_data(1) <= i_DacDataClkLocked_p;
          slv_ip2bus_data(31 downto 8) <= "000000000000000000000000";
          slv_ip2bus_data(4 downto 2) <= v3_DacAMuxSelect_s;
          slv_ip2bus_data(7 downto 5) <= v3_DacBMuxSelect_s;

        when OneHotVector(3,16) =>
          slv_ip2bus_data(0) <= i_PllStatus_p;
          slv_ip2bus_data(1) <= PllFunction_s;
          slv_ip2bus_data(10) <= i_UpdaterBusy_p;
          slv_ip2bus_data(11) <= i_SpiBusy_p;
          slv_ip2bus_data(12) <= SpiReq_s;
          slv_ip2bus_data(13) <= i_SpiGnt_p;
          slv_ip2bus_data(14) <= i_SpiAck_p;
          slv_ip2bus_data(2) <= ClkMuxConfig_s;
          slv_ip2bus_data(3) <= ClkMuxLoad_s;
          slv_ip2bus_data(31 downto 15) <= "00000000000000000";
          slv_ip2bus_data(5 downto 4) <= v2_ClkMuxSin_s;
          slv_ip2bus_data(7 downto 6) <= v2_ClkMuxSout_s;
          slv_ip2bus_data(9 downto 8) <= v2_RSVD1_s;

        when OneHotVector(4,16) =>
          slv_ip2bus_data(31 downto 0) <= iv32_SpiDout_p;

        when OneHotVector(5,16) =>
          slv_ip2bus_data(31 downto 0) <= iv32_SpiDout_p;

        when OneHotVector(6,16) =>
          slv_ip2bus_data(31 downto 0) <= iv32_SpiDout_p;

        when OneHotVector(7,16) =>
          slv_ip2bus_data(31 downto 0) <= iv32_SpiDout_p;

        when OneHotVector(8,16) =>
          slv_ip2bus_data(31 downto 0) <= iv32_SpiDout_p;

        when OneHotVector(9,16) =>
          slv_ip2bus_data(31 downto 0) <= iv32_SpiDout_p;

        when OneHotVector(10,16) =>
          slv_ip2bus_data(31 downto 0) <= iv32_SpiDout_p;

        when OneHotVector(11,16) =>
          slv_ip2bus_data(31 downto 0) <= iv32_SpiDout_p;

        when OneHotVector(12,16) =>
          slv_ip2bus_data(31 downto 0) <= iv32_SpiDout_p;

        when OneHotVector(13,16) =>
          slv_ip2bus_data(10) <= i_AdcPatternError_p;
          slv_ip2bus_data(31 downto 11) <= "000000000000000000000";
          slv_ip2bus_data(4 downto 0) <= v5_AdcIdelayValue_s;
          slv_ip2bus_data(9 downto 5) <= v5_AdcClkIdelayValue_s;

        when OneHotVector(14,16) =>
          slv_ip2bus_data(31 downto 10) <= "0000000000000000000000";
          slv_ip2bus_data(4 downto 0) <= v5_DacIdelayValue_s;
          slv_ip2bus_data(9 downto 5) <= v5_DacClkIdelayValue_s;

        when OneHotVector(15,16) =>
          slv_ip2bus_data(15 downto 0) <= iv16_FreqCntClkCnt_p;
          slv_ip2bus_data(17 downto 16) <= v2_FreqCntClkSel_s;
          slv_ip2bus_data(31 downto 18) <= "00000000000000";
        when others =>
          slv_ip2bus_data <= (others => '0');
      end case;

 end process SLAVE_REG_READ_PROC;

------------------------------------------
-- drive IP to Bus signals
------------------------------------------
IP2Bus_Data  <= slv_ip2bus_data when slv_read_ack = '1' else (others => '0');
IP2Bus_WrAck <= slv_write_ack;
IP2Bus_RdAck <= slv_read_ack;
IP2Bus_Error <= '0';

------------------------------------------
-- Output assignments
------------------------------------------
ov5_TriggerDelay_p <= v5_TriggerDelay_s;
o_CoreResetPulse_p <= CoreResetPulse_s;
ov2_AdcRun_p <= v2_AdcRun_s;
ov2_AdcStart_p <= v2_AdcStart_s;
o_AdcDataFormat_p <= AdcDataFormat_s;
o_AdcSpiReset_p <= AdcSpiReset_s;
o_AdcResetMmcm_p <= AdcResetMmcm_s;
o_DacReset_p <= DacReset_s;
ov3_DacAMuxSelect_p <= v3_DacAMuxSelect_s;
ov3_DacBMuxSelect_p <= v3_DacBMuxSelect_s;
o_PllFunction_p <= PllFunction_s;
o_SpiReq_p <= SpiReq_s;
o_ClkMuxConfig_p <= ClkMuxConfig_s;
o_ClkMuxLoad_p <= ClkMuxLoad_s;
ov2_ClkMuxSin_p <= v2_ClkMuxSin_s;
ov2_ClkMuxSout_p <= v2_ClkMuxSout_s;
ov32_SpiDin_p <= Bus2IP_Data;
ov9_SpiReadaddr_p <= slv_reg_read_sel(12 downto 4);
ov9_SpiWriteaddr_p <= slv_reg_write_sel(12 downto 4);
ov5_AdcIdelayValue_p <= v5_AdcIdelayValue_s;
ov5_AdcClkIdelayValue_p <= v5_AdcClkIdelayValue_s;
ov5_DacIdelayValue_p <= v5_DacIdelayValue_s;
ov5_DacClkIdelayValue_p <= v5_DacClkIdelayValue_s;
ov2_FreqCntClkSel_p <= v2_FreqCntClkSel_s;

end IMP;

