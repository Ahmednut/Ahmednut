XlxV64EB    1871     8d0*&�`�U�ӭ7�g
*��ٶ��f�����ro�㼨LP�(��ɝ�Z7�w����O2h�\��5#�5��L*y��Q{��
0��*�떛�2�l7�n��k��À ��>[ҥ._�z��Q0[o &�/��M��Z��R� $ pI:﹪�d�%V��w��[��I�J>�F�s��r��;�a����wKC^��>�N���'�_��zq%s$��u�s��vk�3l�PkJ�Iu���-wݮ����LO�s,�H�X�k,�|X0������J����kh��'%���o�n�m|TBbԊi����T��~$G{�n|b�oic�����=}�[)�Y���j*��E�|����-����iЊ���u�x���5,~�Ed���MG��FȽz���k���3��(T�-�w�l�g!G?�ݲ��cg���.�T�W�F�A�kP�h�d�`�ڼ[��~�?�i8Y˕m�n��[��z3_�h[ϟ ����z�������-�Z�fն̴�-�	�qm���-�m�KC!W������1�<|r�O6�EDzY��� 'xw1Kr��
!C�g��.�bOs�ݗ�y7�6#Z�j �S9���פ�F�Ei �6Ʈ���6��2���/ �J����f&��i` �qr�^�gN�J���~��l�m�d�l8��" ��E�sXs���b����.S_��Vu�vCxhP�T�ߖc�i���ؐ�9���5CbJ�iY8�]�#X�B��~~K��F#�f0Ѷlk>�S�����Qk��5x��3	����hC��@b	i	��fn��`A�1��E�>:X�hՔ').l�2�	>�yH~��E�U�G�o	�x$�U��}��R�u=[7�\���c'����ya�J��n�v+��y�����7C�)+ö���b�N��^�~>xa�E)�	��#ܳ ���I:��~�,�,Az�㠤�;Ơ$-��P��s�>��m�i,)A'��I������.�S����Ƴ.�wગf�K�A��H��+�@Q��Q|�;�	�P@>��0�EP9�������@��6Vk�2�3�p�T�P�s�/9�8�g<�M�#GQ���8�ge�8>Z�A��t�%+�wsk��xFo�8z�5��5 ���8�3�u>G�K1W�(���8�r�%�'i�X���{D`+�u$���@��Ȥ��⛛z�?,K��F��uD��'�)r�9�N�=�U����Z�ĕ)k�旬�,6F$]t���[Π*;��I5�1��%��gp��(Qȫ��i�t�j��pْH��f��M��|v1�7ܿ�Xh$^͓����Ux�N
k�a�VIͅ?�>خ{�H)щ��6<Ђ�}��`��2ې#E�Mȅg�u���6`<���Fz/�h��5�o���X�a��}�{�����6<E�b���H��b}^7Q��wռlY�>���z6_�u�c��]����$0�(o{)e�}�CbT_�RO`����U+a�&�le�������M�U�5�r~�D�ߚ�7��ǜf}G�_}{ 5�b�n5uf�a��7���=&����ЯGzDn�Z��ڌ� ��0H�n��?�kVf�~�Ҳ�~*�2YY�1z�K0��8�x���))LHm��>��"/鎹j�����<��2W�>����[N��C°�a�8P���^��dN4�g�+
^���3rE#�[��B0\>1��|`�z�����@C��O�D�!z����;C����ix�l��D����G��������D�z8��t�/�ܼ8a�Q���%:��6i->��-�E�o��v���i�4�aZ�U�4�`>��#t�A���!`�W^5�T�MM��m��@�!?��]���?ᑂ~}%�`}��r-ȉ~+A�L��i�{�I�To�z\���ߞxm"HƦ�E��q0���M�5�H��F|R̤k	�����u�b����o\����Ψڎj�HD���d�UW1G��Ca1��i���VԿƌ�#Ğ���d٨�[p�*-`������B����A'�҈�~�P+?� B�rR}�-��D9���@}�xd刿|CS��nj��5l?Utq��g�_�����x�����vg���K��N!S��J�hu�=�Ôs8�߮�H����s��~��n�폹�X_�}2jZ�ꕔl��Q�rMR��[х`�� 0��3H�f}ZA�/�c��k�\��M�%	�����e���J�K