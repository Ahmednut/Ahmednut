XlxV64EB    2e81     cb0��:�܌�G���o��=P�����#2j��^�o��R7�'���1UNgAvXU�fH�L� ��1�7ǋc!>}޷��u�a��J���4�m��p����z�$�y@�/2��X�U(汶"г�8D�G����%���ƍ����@]�Z �4��t�^]<�a�ml�%G��ᥤ�tg񞱀��o����ڜ�k��s����V�3������ʃ*�v�sp��U@�!��R���@�P�j��&���������eN��[S��Nk)�Z-��c̞u��"���ߖsn���euwT/��M{��T��٧��#N^���p!���E�c���S_E � A�X2U�)q��M�:p�BL!i	�i��&��j�B��6VS
�d���𶠝/b	�W�a��kse_[�cѢ��{s������_���]X�6m|����߼�3,���I��ӝ�B��&=��_7?�>���ů��M�b����.�E;�,�����F�Z|̮�C�?��a[���og��h^�B�z���+]���NN�#���'�����
�Ϳ�e&�7	Ƅ\0a���sZ&SgP��qu}��&Ch�q��z:p�M�sSx1V� G�z���`nr�2����,i�"�⃠��M�y.m�=��>J������aݭ Bg	�W��*rU�{���N1��|���vc�=	L���7���рӋU�UT�y;��+K=������Y�t� N����g@�=z
=@^����~5n�����A����/)jn��c�1�[n�@-r��1�5�kg3E��9�E
Y�e��S�\�¿��q�')��|���5�����|G�6[�3�R�O	ؼ�Z/��23}@)�Q,,�uĲƌY&7>����`����Yl�L9�d�2�My���[7p8�;α��X˙�3Ʃc3yi�~G���@�YԔ�;�����g&�_��T�F� ��oQ��G��:W�c��+~�?���k)�@�!����E�I:��O��!�>j�BM��eT���+kI$޴����c�ܓ3��r�g��R�:ӯF��>l�����c��r��� =,˃Z"G�D��������$�M���d{^2��8	D�	!�u����-�&�<h�i��<m�t<�D%UA-�ښ+��?�B<����E����@���L1�w���#�r"�{�j�q<.��	�Kb�c�V�u��ܖS���L:��J��dP��ӣood;�G�SN_i&|q=&�6/�G�dp9;���T��K��K�>(��	���eૻ[��MP��HQ��Y/O�&�����4l&��Ik@��8]�8iXb�ҋ�Еߋ����&M�U�W�0x��*�Ps$�(ԙ�<p�Vn�	U��Ő^w�PAu��?�G[��%zd|�l{Dר.5fQ;[��-�����A� ���z�@Ҍ�L��~�$V�t��^��_~[y�I�\uk��{��9�d4�wE�Sn�'�o�	W���Ψ��/�;уÆmS��*��\�Q�aߨ�czHb�ZF�X�#}�L")��^^R	`+#u�3��sI���l��s�O�w(>m��f�iPP��k^@�i�����������~f�4�o62�Ѹ�he
;SU�SO�:��̭�)���<�pq�j�� ����M#H����應�����U7X/����n�:��� ���$m\dD�pWGR�`#A�?�s
�h��qn�G�I�ΨB���e���p�P��&���m�s�ȳ��o���37��;F�����&/�f��B*b�/�&^���$�=
�'�L��; ��CxZ�R#
���Rè�vT���Q��/��=C�"�ب�V�y�ߊnk�ې�^͞!��3�XL�0���	��-Y8񖙾^aS1)�-�&!��(�!��}ǷOgc��1Uj��H�z��3��*������v���s_�>�6�IW�uI��n�����h�m]C!�z�`j�!���^GP�k}ܔ�!���vG�0��� z��	�刾"���Z�	.�sg�Cp�Ⓦ19q�2۴f�͑ahH}Y��9a!%��p�!��>�7������GO��t<��0,���Д�Q[s�#`Ă��Ӿ$4?�1K�O���&��to�x{do'ZY\�GM0���o�ؠ��0K	���I�j�:�����M��R��5�Ͻ��rS^��t{��/��$"	���a��,^"�f���d��r2��{T	{���)ɓ�=�����Tv�N=� d�4Vj��:Fd	5	��g�8I� Dr>�X'#����%���z3��������
� �.~�(������m�1��Z��*`BO>�)y��(ԗp�2�~�hܻ:j�69��f�����¹$��O�BƯO�����I\��5l2��9�JC@��fm�Ҕ�?�J�5i/y�r���K�Dus%�|	]�|�l�{v�*��TM�)R�:0��/;W��=��G�ļN
�^:xs�ٞ���_�- �L��WgTQ��b�*/d��ЇV�k���f3���.��
C�;��@�{e�&��*��ie��uպAy���{��X��.7h �G�		3-3�k�OW�V�l	��q��-��/y�R�o�����y8`4�6�:ph�2	�h��3g Z,�h ���Bs�s��*��CU}P��W�����?Ec$���$9De���RT''qr���tEJgM�\�;f�SB4�/�.jĖ�*3��׊Ĭm��9��3�e���vq�aTi+n�'�M�o�2��q���=�79�&����"��q��[3���;x�4]��㺙���ZwB}-"�-�Ư�����!ép�����}>�o�&���D�C���,t�K��jo�u����@Ƴ��{ A�
�^j�����obu�=V$��pdv�X9	\�Es�h�`0�3)�}:�<1�~Ih���-��lSqx�ٵn��t���s<���±Z	L��a;K�L}3�0��A|b����X�9 �_xg�v^�6��Tl��,��U�1��٫X]1v�nmxth�<�M;yJ�Z��c$���{�d�Z?]�������ژ(���Imn�t�[�>!ԋ2���g�0��S����qu`X�|!���l6x��)K���*y��Ͷ�aV�)VC�*�k��-`u�E$(/r�:1"V�|��yS����Z����7aC���:�
�3�y�6�-r
Xp��G��5_���Ԑ���:��{�