XlxV64EB    70fb    17205jv<�_A�ҬO�pQ�2jH[Ĉ�+t�i�5��P�#ـX��������y%/<鋷*iքD���ʍ�;�7��~)�y�~��������n��$Ó�����D!��/pB�C��줟��-�a��2A"M�;]�M�pP�>"�ʟj�>�2�-@��v#�*1��G
�����?�DE�[�װqz_І$�FM�UH��aKR���	x=!��$}׀=A/U�P&Z���D��ݘ=�X/���
¿+��3��p�TS��7}NrŶ٥Ⱥ���^����ݯM�������t,�P��S\�}
 )`5?�/�^I/��!���{_���*R#����+��A�O��2Kz~x�
���g����e��>��ǟ�fN���eR����9����MPش���S��%�H��'���ؗ�C�KZ�� l����t���<
s[J��Vn_#���3�V(��h"��(~j�P� ��xb�&��E�wR��m�B�PF=��`	��Gc˺
�h���[{��l3�ءo9.�����cU��Y�'!!\v�u1Y'��X�m-���y�~,�?e�\ڷ<�K�Eq��b�͚�ނ�xކ�r���ə�P����;�X��h���(R���	�Ñ� f�s|���<�J�}wRj_?}�Fum���$$����[��S��Q�
��vXP:l2#ϴ��<tX��IyN�ԭ�*�n����=ΧP��BŒ��mGC�@��U&¶����1�P���#���F������U��~86�e\ �}N���8����^`��4��V�'���\�ȍ�kBn��(���
��"�iwd'L��j񪿝c��
���=��S?�ft���%���7��m�Y��b���U�}���ٖy�1��j���=���#Z�@������N{�l�6���P�/|��
s��b7,��T�-�Lq�6)97��+��#���H�$�5����h��k �2W�б9�b�F�.��ɮ�$�	���=��9D�~v˷F$`��� 'L_��g��`�J��/dO:����:��u��|��6�I�����b,A�E�',�g�AMFc?=�*q���NZh��=�G~�?�����<�y%Z��aDrvn�AG07Ƿ���ax�#㓵,�bn�|QZ/)JU���ؠ�ѥR؃��(�	!�I)�W%��,�!���3�C�G���6�ٞ9Tl��R�^���Fݫ���/�WBF���Tiп%�q��B7;�$��
 ��*�/RO�T�g��Nd,k�w�R�x������x!�L�DQsؗ |0uQ�a|R!�p�� G��*��#ҿd
�>�.������#3�@ ن��:c�#@+4����}`���j(|^�����_�O~�g/ǈ�Ю낅��RLu,.�h��hB��m:"<֮�U"TL�ŕk5�2Ia�ϋ�^��gn\#�^@�e���
�e��@PG�'��w5;Ɋ[a�& �'\���BUx�׭%߸�tf��Z����ϰ�a맠1[�x/b��a:�'S1�ƶ�`�<W���г��v�kml��P�ts�i^����Ey�Ϝj�6d|��]�������N+H��L_��1�(ʶ�뭼K�}?fqӒa�e��J�[d�ѓ/��w�:��7�J��X�/&Kr&.L��̳c�������J�9�S����j>�*r-�9y���#�.y�������A��^�S�������~���_���0W���l�������U�ZT��0��a���������X#���O��,�*>��Ʊn�L(f�m�w<ha�e��IO\*���W��.ύ ���� P�Ѱ ��ڵ)�@I,nF��!�j���VHQ�(Z?)�y�L�""�G��(֙���#�:�`�[�6��f�-��ڭ3�JF�Ll�ȅ���Ƚd���b�l	�g���{s�&��ʹ����~C�3��w�^B��Ūl���CȞ0�Çr����C��vH@䗢�G�ѱH���+�Z'v�ږ�"�黳O�g">�?�~Í����8>mp1��/�ÿ�/�1���8`��f���B�[T�v�G9]���s��2��A�Ϻx2��_"v���}NE�B9��	�YYUy�u��T���+��9{d=�����&����\�b<�nG'�3k~�9�����O��M	�*&k��R�2
�E��V���X��0S�/�	>.:��@�t�������B�l���*��(�U�ސ頲m�3�KS/�q@�&mU/g*�H�X�y����٤å���������/Uu��b��w����l�Q>�E���� �k�^;W�즧��6�!���a\��3a�_��v7	*�0;�9�P��:b��љ�neMFt�c��m�#�#��ݦ���zft�Տ��������F�bDh��"�r�������;s��]�*-T��1�֕�
�@��2/Ea/z�Oo-��c����7�ƑC�9^��bA%bJ+Lł�tP��ցy�Ϳ�L^�����A��>�����B�E��7���~�2!fn?9.��@"��2ցd��+�1�����65Q4)�r=z�����Ӽ$wF��-8�1ȹ�/�T�oA�/�F	pc�!L�Ni�����S�x�� w����ݛ�I��Zqe36�Q��a�COKMY���\�}����n�H� Si`7�*�Q`dw7i�I�?�O3'%�Bg���.PT.�3+��C�d�bI}���v��H]Avs������5�%Z�B�"�.�U��g�]z���«�M�j���
��g�$�&�Q�ߥ��	,�θLN!�Ȫ��yЛk tm �������Ed�S`�)m�N����Ą��8[3����n$'[ߘ݁F�'"A=��Ohi~�-�~C8D�=�.J{�t%ӫ����1]\��H���^��8LvV��iީ}Eq���0��3��c�,���	_�?�ƕq#x�ٰ9����kD���W8�aZ�59���n�����d<.Z�%O���ӘW଼�AU�cj$d�nm:>�2̞�U]�T�nE�Pgt�<�9>����o�Ii!���X��t�8��6pM���p,���g_�NV,����U�bW�Ԃ�(��
���e*뀕�:�eJ���F�Qv�+{��0�_��]�.���9��F�n��iG��̢�_a��9r�>�/�0��3J��	[�_iRK�վ��x��d����u���� ?��������$9U�<���� U\8�|	�.dV�
��6�Y��N[��B#:�Gj�y���6z9u( M��R�IgܚP�E���D<݃��V���m5��c��PHW�������G�2�s�d���!\@�`�O��I��E�t���gZG�>��ܷ�HҁX��N�U��= G��`�x<�]��'�`7�G�VmP@��'�4	�"Չ�i$�e�tH�'d�_(�����-P�f��W��Y={Xk̦�у���8��uȒ�؛I�(���̃
�J�ݗ����N']�kMJW!��TX���N?�����s�v�KzUכx���c��cDS܎ ���e:�BG,[^Ԛ[��ZR�_W����8{�Z��}肽�����]��4ȂJ��1���saOc1�v�C��,�S�کܿ�Z�H�4쪭{��	U���^8���{��3P�:��Q���p��6��x�h��G[1rW�{�Q��Nl˔�I���*V)9��gМp�U:#�Q:פ�۟�>�RRع)�m�|$��ɾN5�Ds��?N}K�����z�ck�#��^�����`���1��{�5�TC�;7A�����Nj"�)����{(�(q]ޛ�ux�i�-_���,o�_H�K�B"v���� v��\��AΗ�b�l���(c��)�-ј.f����3�^�Ph��h_(��g>�<�o�Sͯ�i~��}�J��1AT.�<&�w�
�JJ��9�h-V^)�&�(?�
5�[-̓5�vFi���yi��#ώ�5u_i�uP`���y�e�����e|L-������x�S*'� ��>|S@��ʍ����ҵz�E�Z!�u#1i#�f���]s�ve&䆷�����'w9�ʅR���t�:��Dc�[ӬN��I��3�G}�-ࢽ6%X���9@73417��𬐠�6�����1{��2���,�JPu����NO;eY��*��d���o�,ZP���wzm��O��	A�%MYy��k4ɟ��3<����O]�p�xk7E�|vӶ9�E��Q~�O�_b�_�|P�� 	:A���ms>{�1�r*Εd�XH��cZuL�T�^��SA]Ty���;�p2[b�z(������nE����?d���)��n�L�ks	���gV�% VP�����.�0y���Lېv�.z=�E����}1;�[�X.�j�^�V�f.[S�<d=�^p�{\�[�b��̿ב�#���B��y]��D��G;�{����K����9��"�ow���U���A�s�4G5�<�U�4����>[鷠���gW����˹��69r\I����՜�%}G��ME���� L3�����`��iyzy��IG�0}��iC�n;A�2���M�1G����ڐj0��J�y��r3#���/4�BV�N��[yJi��8
�ȳ�n�U_��f�j\N+�Y����!_ ��ʲH�җ�rmu�f��(��2n7n��
ڠ����V��X�*ږ��_
7����6�p�qmm�V�����k$�j���H��bJQ���0��2�B�2#��A:����`�NY<F/�4�Nf�S���H��fKȋ�)��\=_��@77v:������*�����pR5��ؐ���W�ZeYyky��@F5�x����ά<�������Q���S��8A}��UM΂���a,J�P�5͜YB^���=�դ�kZ\�í@JBۡ�����ǀf���9h���ͬO\8�����Ӌ�xh˵��Z�߽����R<?��i�����D]�C�$��S��AoXy&��l�6Zl�VM �M��3�����O�u�Q��')��h_n�ؘ�����]F������^t��l?P�e�k���}��+�0���N��b��<ys굦l��4j�:�N-9�K�ߣ�k_�mC��e��Sk�D������I���E�8�9��C�1��s�h�)��%|���� eܜ�rN�����2�wGZ�8$S�����L����n;��uq����O�t�unǰ3Ut=�%���Tf3����9u��Rǲ�_&�˜;	
�~{X�> �Oe���*h�����U��(���P�'�^T(���R��BDʁ]e�?y�}s$'��2U����B���8D�����j��-C�}.�U�F4Z�>:#��1]��@���N�O�b�w؍mi�����R�(�l�>���Y���9+�c���;'?��1�:�+�6�I�-��R�LYU�9.�4G�������e�Yh�غa�$0n�o�g�)"�`u��Aq��J���v]�rp��^���_3iz�?��1�#k��)��\0�Μ�\���ӻ�R½�#ٖ(����B��
����c�}�{d�����D4Yb����~2�%���fHi�UPǽ��e���� �[i}��b,ʨ��/B>|����X���0Ü��i�{�!.P5T���Fm�ڜ�rlj��g�W� ��lj5P��Q�y���(�#�7�Q�|_���%�sx�/�O_���2���/�����q�l]�-�