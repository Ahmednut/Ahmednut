XlxV64EB    c849    2590k�S���4r=�xsϺ-�r@me�l���&�����d�F�ɕ�CO!
H�_+��h̳a~�7&	�'x��t��K]���U04b�|L2(������C�����b`�C��Mgm��3L��I��#�ȭ\.���$`���~b7ګ2�5E������(�J�8v��7�f݉5]˭o�Zx�ܢm:^�j$;�0^����_���b]��
��id�0���C��"} *�����Ĳ&f\Ү���%�B|\��K�l�]s� �h/d�޹l�*N���*%�RYo���9�.غF�Z��L�|�}�m�ʠ�%���7���$(����񄢱ݕub���4�4�k�;��iA\��2U���*:��u,p�d��zy���(�^g}2V��M{�
�p��Z��V� �y9g�+�IX*O���j*�����+��ֻ��:ٺ�WZ'�Ӓ&�fU=�qY�)8�j7���� u�H$Mk�[d��.��fVL1) ��,\��ӊ:��(��#/�
��(͂~��e��E��,�R��O�
��<��5��,;�<^�_,��ܛ�崧]�Ƞ���0�΋��+T�4����Kgp�x���Z�p;�8C/�f[UQq�j���۝�I5
�{{l�[�2�薲\P���Ȧ̞�x��Q���%��A��ߊ��� �������� ]#�N�Ю�g6���{H����PZ:����G�+���s'�1�	�j��$g����8���L`�}����n�&u;,��no��FZ��(mh\��j�dP�0��
��?73�m=�mS�^O���Oċ��8Y�go�uA�k|LA��J�q��"�6�C]�4)�dZh��#�-�'����O��%�s�!�B�
�}�S�no�вK8c�Q��[Fɰ��F��kE���ձ��b'�@� qk���׿>#h��ٺk�L�VoСF�r+��a�B���yU��^�w�Y�����HL���t�B-|��XA�/v����YY���+�
�-���&���H��|bw��.V�ln�h�7�䥯�T���^����=��b)�B�E�g�Ey�
U��h�t��/aX����rCxX�*�Z������J�����r�6(n?����Ǔx`X׍��|y[�E�5.��Ul��<�ݨ(^6�jo�l����G����dm"9+�p�h2󂥋��`d�<�h�M�������ta�H��m!�c��6�֠���9��wBn������i�9f�4?���������DbF�86��d�Z�n��yE����d���i�(��XX�8�kojhx6n��H�_������vJ\|$�ܷ�@ob<A̧���5�nن�E:]�^��zm[���0�yX�3fh>ci>�-���?\���3��M�csv)[Q�GU�u��(E"��J�ڲ�߾Tu镬�ݣ�,�b#�&6!�\������W���5X5��UU�K
}��.룶�.�'���j?.�#mc��F<C��H�|o��)��Z*�`��)A���=�l���6��� �3�(�a��X�r9B�ĆДnsI�Nf&�v�$�)B���T+���P~:���/̻Fc9i��+�Mo����Ӝ�YZ2$�A�n�Ie�N8�k[�$[�3z�ʫ�;��;�sM�[UJB8�{�ybv��JF����Xr�jH��j�.�4��ߡ��F�����l���|�o��u�>�y�/)���m�5�g�SK;uۮ0t���ur�2 L?�
��B�l��3׾>�%_�!##F�L��k��0����3�"�S���; �S%�@6¼#xlC�}q1�� �b��&���n�N��[���,����r��5ߋ�%�6��^�c������7�	�b�%8m�n�������]���ݿ I"�Eoon�)�)�����4��x(���������M���e]J��l1:�(<Q�^RsIY?���s��ٰ�tA���9�z!.�>�wph���\�}�;,h�������@G9�Vg�\��M.{h׳D�O2�˿���QQ�c�lW�jt�g���^����+�)H�1ݜ�F��E���YK��?љr��G��*&�Ba�6V�����98�zT�U�0O$Ҝ]����I�ْW��]�����h�e��z�#��bdX�@��;[}�@ơ��gS�����TX�0��9�d�j� �(L3f7�vЀ��Z�Z
t1��{���-��'Sz��ݽ�H��,�S�U޽9��i�2�a����:կ����q�X@rV���Ek;nW
+e6K�i��gV����ue��9��,��� ��:`��iE��H"l_��"r4�9p&�]Z�W��������ʽ��l��j�`t�'�0��h/�2V�k~kB�y���_ץ'U�/`l�=vРD�0c�{	��D_G�׷H˸ߌr(�h�] �Y_����C��)k,��Pl��uq3�����T�G9g��E��l"X\V��'y��A��ХP���ֵ�u?��|�uЍ�c�U��!0Y:�QEJ�(S��s_G�]T�u5�M�s��\������d�IK��.58�E��-��Jt)�,l�.�IQ�1��B2��lFFn0ۗ�ݞ���7�i���i�@�ٖ��=cB���=VK��T<�܀�y~\�Y8�ГI2���?/�:	��v�ɟu7Ұ�U��pA������mpBv�EI���T\��"/������,d�H�C!9j:�JJh�"f-L�h��"����}�i:����(a�ė����>�O$�uץ���Uȧy�Pp�T��,�i��k!�oviC&�w�-'����X�������ޜ	(���hو�b����?�Ta�#�����l�U�k�5B)O:�8�lB0���z�+)y���ɲ9��R|�G%X],9y��ub�	=��wH�?�@�0�L����=GS���0��7:��]f��S<�ʾ�:;�_c��^��p�3Ձ�m@��6Y��f�����..�}J���=���bկ�j@`^<�r;/�.���d�ނ� +!���v��&���<l8���:��lj�Aτ�$kξ���Y`���V��ZH������l<�(u��:�ː��oi�8�8�ě�c�鸁�x����E�,�D��/�C�+ww�UK���jQG��U����9I���bh�NU92���OGG������b-���f�^��[���ե�jv��P�k�EM��T�-��o�l���F��
��V������`�������5��T��3����w@��"pWRN��OnU6 ��+����Y/8^2��/����� T9s�����n<6Bb�MmPb�b�VAT�B���m�vY��>���Jt�������(��O�bq6O�y���x{z:���z>�Oo�w@o�V�"��b�B�ta����n���pB��N��p�\��G{^h`4�$V'��$~V���;��m��~Q��*dAύt����je�0=�q�����݂�l�+�ײ6��۵k+U���9�,a��|��޾M:��cOd(W�5~)���*�������_���f����`�H/7)_v�����A��b�£����J㏻�Jj^�����$M��������[xp�ѮL�<#'�p���7 v�dF�ȭ�Mt25P(���C�����2A�ws��c���T�T�t߫/4Ak_&����%���B����F���5���6��]F�c�� ����yȎ�u�C���,k��k�ڽ�X�[z��73t:��@#g�i�9�!�/��-Ï�bNY�]�&�(��Nz��r������^�ܛ<�.�HD=V��;vt���*�>鵧xܦz���&Q�4��s�!�K���� ��sG� չ�Ѷy�,4�پ�=��K,RV�ۡ���x�h�l�8��`���V�8��e%;�D�N��q�m���5e�w&��`����~(1��W~i��7`��R�v,��k�᷾#���p��t󥢷��՟����.�=#Ş�%���4� �E;���5��;�O9~��I���ғ|�
�^�o�f��d� ��.K�N�R����� ܃:�[�G��Wc�.�M�ġW��C ��*Wk^�\�� �;������󡦎�Wڽ�f��?���s]v�=�X/lR�[\�k��R+g�K����dd���Oz�X��y'tШA�j��&!���~4�R�U9zog��V�19�P������p����]U�т��c���<(nbOǯ�oS�s�{S��.���,�̼D#bk��2=���p�_���z�|��/�,�D_Mt̳��5�p��@/҂:C\�Z��(�	
� �k0�RW����'6|�]�Zw���<;|��7�m�|g�"��S����ҝ��w_��c�@�)h���k�k��ݡA�U!�������
AD�~Q���J'/ ���ӎ�j�K���å�`�RY�;4���2PI���k�����5{�1�aKiO�O���3ױN�V2D�n��m�ң�'_��I��V����Mֶ����2
�Zגd�w�D��#�kSv�R`|D�򽇚�0!f�����o��?��2P�O�S.��]xu���"F�H�%5�?������Oh|9� ����w\]��\���&Z!��vRw3����s\��z�h\j/<.��u�I��c�W��2�ׂ���V�����������u2>�k�U|� �sx�.��i=���/����qd�b���tif�eӦ���bԯ���#5��Lp\���%��M��/mCe���z[ѣIW�q�Ju5��
�d�(T?�������R��*�o��;��?FYQsd��K�J&�q��2n�b�yk˕Q�m�\>�\��`��Y(0h)=��5�h��;����G�#K`Y�y�sOwٶ[�2NBO �{�N��߄���i��6���a���K��~r���~���5Y�2��rď<���[Z�^�&F��h�yn$���˘�㸞qFd�J�[?�cY#����Lfu�xM�0�t,iA�{���7ƞ��csn�.qM~���a��Y©l���&���x.Ǜ�*���Hj���v��D1�#HǴ��{s8>�г�y��7�5ak���#F{#)�;�VrSA\��?�N}tw���G��H�{����]�B9dX��w�6ز�&��ҫVL��9q��P�����oqK�'#���k��&?�T���$F2�fq� g�pVG��i�[d�����?�"�U�8��Ǣ����ׇ���/|��Y�\O0���]MS-��������Nu�#��E���]�D úrT;5�W���e��q:�byЍQ}V��UxM��3�̟�Ai����s7|+��!b��J�e>+��$uR����EV��i<woR��:7}E;�%�]+�0k�P�ؔ�����5�<2�r,�A�xb*L]�m�U��*�k�u^�e|�*��)e$�ERK�C�{�*m��g���s��*�\���~�V�g��ߪd��-� м���'�z��M�`\tq\5]O"���4Fr�x����t��4<�:���� NU �C�dݪU�m^S����������洙�!��R�2�xXj�s�=�|h8���N�G�X��c	պ[f��qr{/QBr�T�!8{Z�*X���6¬�<���J�b�<^�� ��PXw4)/���v�|�[�mׇ۾:mA���e�5��ǀ�d��ٹ�/�bŜ[&7I��|�,��5f�Ϣ�]ݚ<��r���+�9��i_��!(0�1%I{	M������ɘ�_�V�+
��,��9/��.�G:0AIc��^�In_(��+:sՖ�=�O~f�#\��f�#��?Ԇ�A���)C�p���W׳�(�Jd������	ؒ�ۢ.�h�F��Q���@&n@�o���6�DA�c;7���xź)z{�Åa"�ئT����=
q��������y�;4|Ջ?��W������d��B _t�1}&p�?�oi?��.�`�\p�@���<N�	,5��&G�?�F%<�·_ŇlR��D�g�'yDp�0>|�i��&�D��� �ޠ��+���=���"zf�7��sa`����4���L@��+�7Aaj<��A��SԚ�&U�o�J�%�RG��B�9M6\���Y��/<d�W�Í�����01MO(��gQ!ڇ�a@^���Y:�?F�,��Gb� :��$D��M��/��G�7�g�>�ʛĥ�����V�l��S���<�g\��\u#�,Nm(�ϱoDYᵞ3Y67�I�_`Z�?�ǡ�x���ɞ���M��sl��E{~�П�N��da>9�p��9�)/"��d s�g�|����|�U�{��g��U�p��I�Ѱ�[�cM�ց|�<� !��_F`���C��[�u;T�M�:���P�u$$Ԧ3
��тȺ]��˓��R*9o�K�]m8K���_HN�"Y)X!6�Hǟvږ����9�B䇺�e���{��
�{�<��q_���X_�Vl�*q��[��ޫ��`��`������Yn5y�TY�ڟ�@L���(z��=`c7J2�{�FUxD��Ћܫ��3v���vSqF����i��O�N��x�𰪧A�8L���׀$�9��Ǿ)M&�B�T�D��-��%+�z?��k��~M�j��7�R��F�Yr�sɐ��w8��,yk����_��rU��xU�w�Oh�1�Z¬BJJ�J	�����kTC�D�O%�)E�<bgʁ�����T����Ms�E���^��2�=��l��D��b�h�d�{i�,6�D~�2�?��^/�� BR%2�ӷzW����\�2v��d&-�DÜ�'>�q��Q+^��$��tx������@��u��������Dz�T��Y�y��S���ԽYu�W
F-��������d赡�g�S�Ќ�6"/� N�A��xy���Gxl�<�7wQE-l�}+Pi��2�^Ԫ�ƻC6��~�(��(>6���"����n��@�%F�\@�Ӈ�S�W-l��pD<�Jxv�k���
=����`����Go��Spp�[���>IJ���3tc��'��P���-�����,K:�C�[�������ߙ8���%�C��q+���:(����mڍ�k�/q��E5���Q//��w�ױj�Q�M�gd̖d0|,3�@�[ݚ(9���*�a<�E%�=!;��Y�;� tn[!��o+'�J@��]�?���TF�?\;=��(X ��|4��%��E"$!�����J��t�F�)z+HP�pa������-��~����c_��o���[v��P��
7h{,�����>{^�%6a�L``0,���=H$��^=��_u����a��r�ɼ6,���UW�L�՜�����♪�����>��f���nj�l�c�/�Oi�:s���fB���u�MMm�X�J�K�A�ģ�5dG��k,3ͷ�8�.��تf��=�1�����2*	~���g�@Q-�'T�����{�h*O��/�L�Ϻ�����w1p��z~`���_�����s��1]k�e�vj�����o �fQq+��e��bJ��E�:�M����p��<4m��\i\L�����{��^%�d?��1�Kp���s�V[�X�a�.a�O!?=�?���&�<lcY�h��s��v`zo-��h
������43��V��&������k��:�|H��\OoW���ӷ'�	���o
)@^~�Bٟ����U�Hfa��5TD&.Z�O�s�ݖ�<-@�ek�։%�bP�D �=���@XdݜI���*'�=��S�%މ�~��X:p����(�]=ի��)`K �K�vms&�'Y�;��ڼ+�$��ݸl��w,`���X��M�Ff%65nѬ�(Jĸ�jF��T�Z)fZ�����2����]�Q�ۃ��6�jk��|,8���q*H��K���P�9=�؜�K��b��?l��o�j�P����q��.76}��1�y82c���W8�I�9�_
x�C�ȉ)�
�OK��;��h��#9��x#5x8��E�h�eïM��^<�stJȒ^ �m�"��Q��N�p�|���ѕ��$�u�#��..�q#SC*y��Y�jd���A�3�0�R�Bd0A��]4�qP+*�9�	s$0=���eSB
����O,�1'��<)=��)���f�)l	=�$��b"��#P�@��2C�_���W�a H�'�+M����k�"�H�i�� _]�z�[%o��)V*{.�I��l��ȻJ�^�2N��)@�C
�$�i����%�ծ�ե�$�x�7L�	��l���D���/�K���b�2�Kf��T����[Q-Ḙi{[��*�ی��!ů?�ƪX��ᩡ���_�?|M��oL���a��
���b~�J,�TB4\<���������u4�	.ޕ��m\���r� R]�2b�U��OM%�vُ�t-��yւ=�B�;��@,n�1��<�*i��w?�\i��&�)�_�����S��M����Ww��NV��c=�F�~/��0��ش�����͓$,/�([�0�Ӧ��y4+���F��hݰHy���g@�e�9%��5�O%~���R��9���U�
><��,k�G�v�C�*��Mk��A�af*#����2M�"�%��Jt���#z���2£p"�`�|�4��'�5;�n��K(�&mzx��w�E���_W���V�'��4�x������̓�%��)�6�VF�"���� tБ9BS�+�
��	[��w����e���􄩠?8��.������C�b�s��e>�1�q��0�_j�Y��Ti;��7,hwv���o�uB���_�d�qg��p�~��`HAqk�Ga8V|V�;���
E�R(7w �<��x��wJ��&<fFJ�0�����ˢ�pS�6��o�F$�LrǐM&�f�5���An"��n'���୰�`r������B�#�\ֹ�������k���y_!�5��6%�H;���$A,80�IGx���W��]��8��R�S1���ɰE��F�8K�c ��N�'�i<y[$!F!�V��Em�n�Qː&a�O�w��I�H{�Td�z��}Y͇8Z�]Y��:�"|8.�垉�WlEJ|�Q/?���X3l��(ZѾOcVͯUn�}�M@�.��2y̝�1�"4ZL����nٷ+Nu��/��%H�t��C��Crz٬O�cv)���%?޾O˽%1\���!܊���S���D�C���sWc�x��H�(L� �:��u�6ՋA�S��\�ѹP%�u~�Ջa{�E|��Ғ%��uk*��leIi���
�V%1������Z� ?�z�/�@M���mW#g���$i:`�vv���֖�q����y�U�K@UI������Ǟ*�J�����S�(!��1٥��J�~���Ʊ