XlxV64EB    1f87     ab0��X:Q�t������u���,��z��r��q���>u�t{��d��v� �-_9ʫ��#7���[�^�E�nD�G�ŧ��LL<�n�͒���c[��5?�"��
r�9~�x|u �,	�e��-`��	��h
~1H�Z���qIDS�u��Uڪ�'�fv�W��+& 6�UYZ�</�������MW�\��)6�T���-�p]K����	Пkt�ӹ��^��璧]�*����������
� ?iM����W�?\\�E�5��6�I�S��^��{.�)fu4�Eȕ����6C	�l��c���)�r����}W��睬�C듇�|�׵��:��I%��ZP/�Z!e|O��$�5ܦ�&�Q�oY�ݯ?ǹ�b���riA��\�EQƩd�S�b��sq�0	?��d�'�W�t��v�ơ�@@Lf��y���`͋���-V��t�"��Qp%@-g~[��JI��,�i~��D�(8�N����e��l"D�
��̄��]�9*�򸿱d{��/�]�����_b���v��KY�ILŔ�/����Ո�?@X����h��YA��X0jT���(1y^"!o�
</Zc���[�v%���:��~�O�� ��?�#���O�C�n���֐ A_�*1#?U?�]+o���{A��Y�]�i�o4+�n�7W�����Uj��N��uqi:L�<ç���fnk���̫��(���@��R���Tz<�B��*ȏ'm��jt���O�4����$�QR�	���ga�6��X�r�v��!�)�9��WΊ�-���w=��1"D����\�se9QbM[�B
��<��j/��O�qѝ����`R����,@qn��L�$z��.d6@�(b-$br5Rb$��d����sߕ�W���"�M,Q��QSX��ԧ�\�M��)�::S�i�XD�Gy)���h��Wp�������.��v�P��t����\��v�mj�0p���M��A�Hާ[(�_��m��7V|5%���W��㻖K45�Z 8�$�HPIW�u��ȑ������DC����)�&\M�1�C��VN�Q��l4�'ޝA��qð�������f�xޮ�Kj���W�i�,O�j8�<'�_�Em��xE�Q��[���婔R�J�H�D������qnP�#k�����Cgn*�?��~5>cKI�-�h%�����u�� �^Eɝ�/��ud��y���k�����no�r���#��� /R~��Fy?K�D >�8��;�ŋ��O��%T�mv����pb�-�s���ѹ�� �B�Hĵ�p bUE���*d�uM���c|r&*�b(�`Wa��Nɷ�'�����YI��zuV���]M��S�2zNm^~�R���"�����q�i�k��Sj�#�[_��^싼�t��=��,n�I����ٿ7��(`|l��W�Ռ����&áH>�4C��{�;�����L|����Ycw���KRJp��d5!������VB��	��ͤ�ʻ!�p��}kӐ�7P�t��@�/�v���i2�s]���6�����Z��5��r5D�r�Z�>��bhv��h�3�t�\�6FJ���K�+���F^~t�M��X9��z�h2K��P`4|�GM�@��P-�#0k_c<��b�Zx�0Dа�/��$�y�C�L��qWY�)*������h#���1�ѣbO$��S�qXp�� n�0�� O�eC830�TC�f��J������9�6�����A��r���Z����B�������"G�3�d�ah! �|ޫZ�g$������ڍ��sg��� �?R������]p� 5��qW�����L�E�^p��`su<-^�j��O��/�3	���s��vqC������Ϧ ��25�_ʀ�̡�W�	�;%���9 ��dYnu�S�a�[��j�#����h��'i�5�0���K��U�H��#ٕ���5O����o��4oKrC�cDRv���
�O��!�Vi�,ɬO�F�ޔ*�B��3�b��jĊ,?�,�V[���M̝`	I4�@�]�!/�&(Mލ�i!⫲���L0��ȥ]V�R�N�
��|�m�˕�n��0�ޣ�U�ɾ��@�֪kr�a}OU�Þ�O ]��}����	��)�k ��O 6'a���\7�jѴ�f��sT��x�ƺ�/�1�^�A�����ŵ?��
���s���@�g�i��%MZ5��L 	2lQ��1��&��GX��X�w��� N1��i�m�������� �e���F���X7A	�6H�I�-��Ô�}9G*�|��H���"�D��U�ҡʥH�����9! �{���f�`�w�q�a�3BV��1�����2�ֶ��r�R�7x��M;���V��p�o'ǫ�R�@� ��c��g�9@�~1�9a�� $�YH�� ���?ް��հ�b��Y�'�����Qb\��`J{�/_�[@�U��E��v�ۘ�+��v�w%�=�0������Ӆ��N���hZ��@I���7��e|I+v����8���p[H|'��$[ȟg�Z���ʤ��~�:�����p�L�!5��$C�on�M��Ԧ3ԙ� �y��H}/L/�tb�]X��G�