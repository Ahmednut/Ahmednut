XlxV64EB    1681     8b0�q��ed�˺���/���:��ќqŊk'V��a)�W�-h�钧E�b��� ��M����EjA������O,r#bq3(�RY+�_�H���~XVq�W3�Z�+T(〩y$�7�ۏ)_M�o1Wb�9�r���,�T"���ϙ���3�����Hag�1�
@}��U���V�(9��5��4Ph,�)l7�N�� �t��u�^�k�!��X9~�\��vH�/�?�p��ẟ��� eG�[$�r�lͨ�W��G-�_\���X�����˽�����)F?��T���sx�n�/���61%��c%���R����
���ߔ$����/�:�kQrj�4�a�u���)�4ӢVVʋ�}UE�3f\d�A�@?�d���#������#bH��l���S�=��n�0Q^��h���:��Q�;vw�ǈ��&�g�u����D��'���>6���z��yR��5M��>J����V����znU�r�
5k���y��W���ړA�؀g5��T�u`�~jGB��/��[��0b4$��w����]�g1$�n�#3f�d3������ً��ʩxJ.���DZ|[������$肏ll�F�6�$�R��,=�$�V������ �F~�O���	�	�i��$._G��um�J�Zn^ �SU�m:�`*O�.���-J�z{�����w�*���nM���[����$%���!�u�w(�y���J�_��]
��n�9�+�e`>;w�<f0��,2$�\n�����@w~V�IO�hh�7r,��a��&�X��-�Js��ݳ����n���&�v�A�q@�w�d��"j������cS\Z��XȡY;$虻lB-|l��ِ�A>w$QHH�g�?ɽWr�G��}^���v7�i��p����ަI�n ��xL�&�������v���On��L��"��A��%�'{���`%��[$�r�_c"9]p�6$�*������s�dI�g�vL��?�uV���d�����ղ�W;��_� �pӛ�GH��g��l��l����ؗ� <��F2���h>�-	y�l�	�o�z�\Lo٨^�	  �J^�J 9�T(N��T�ҵUC���Cm�BQ�4��:r�T����S>�~;�6$9�{�ϙ��|���M�]�����P��� i�!ҿ�����a����}�+uG(gn_3����\}t���b0�a�Ҕ�ٷ��t��\��f��ϢUjs�k���r/B�}���E�����������kT���E|0���~맽�'�uE"��J�֫�x>3�te����D���ar$��@����˒�3s�ݠ6u>2��H�jȫE�� �2,�/B���C#�����<�����sȌR|�nd5��5m�s\�:]�Ń�f'�g�0��Հ`��q�o��+rK���R��VZ䋷���&��Su�H0��i�$E־�hn��|7����W��:��2��]r\_L_��~���/��p �%i)���]��+K�_<��L��7W�u�V�3аlթ�E�ѯg���d{��ژJ��Ҿ�l&T��i����6���Sḑ �v,*�Gb�k(a��a���'yv�E6�x�X�M�,�C�$���H���>��|����J�-.��G�${���`�Vp��wQ��
�:[�V��o�
:X
�k���^�;�3���X��@,�F=�^xB��[zn%~��ѵ����^d��7;U)	�x^��s�lz�N��PC�)�TMtZ��B������fiT��e8��|�+x~�t�~�3��RU�8��۰��p� EJ��t�~I�A���X�Ġ��s�q����̀��7��@j��5�ARƧ�7����^*&[P�� +BU�m�N�S+0ݳ�˫73������=���Ἦ��fU>o���k��c�'*G��=u?���S�B������=7h	���x,*���y��]y
~�W�g�dp�N�/�'$	��Y&�?��T���8ٿ.xX,yK����g����Z��b	fb$���8�C�9	{�tw�4�O�-n�����-s�K�x5�\�mt<=�3l�j���o��lH0��F��J $�^f�.��g�����s(Lq��-ˑ��8�Y����=Չ-kC!SĶ3I	�ˮ��{S��{�߁�\� ����v����)L�