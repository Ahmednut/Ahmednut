XlxV64EB    b72f    1bd0{���8rs�M��2�C�]z�oh4���u	�SrXf��7��dO|�� �;%�ciN�Nc�h�K:�G�xg<�A���
�}lɂC��@@�����i�<��qDK�A��wF7���'�fE�x/�O+ie�goR�m�𥉉�,]zwN�&>b��X9�u�:�)˺����CN���?I8э��Yb�J�M���X(7C�g�ZW��[�m�RY�g鎶�I����B�{�l�6?*�L���� 5{�h��aED�%��U���W����u)��mQ�1
l��:���Zm�����J�[��Q��Q�]Ki��r7zD�Z2���"D�j'~2��<	��rF|"]����Cv
�~F��B�:U��ۢ1�m��U��+�k/���t�;����Y?��x�� '{Z�5�R"B�bz�ڹ^<�F���E}(�t�*f� ����_z��xʏ#Nͮ(��dic�f,�ZGw�ȇe���V��#!*"�W�$G5|,ޝ��pX�`)R�CĬC��o����jcPrC�3������x(�.fD��n���"��C�}\(�4^Y�7B-��
�(�ȼO�]A����)3%s!T�~2�YB���j�3g9��گ/�+�x��uXO�96~�%[E.k��O�|�L�@�lt�F*ԋ_A��K�"'TF=U\��Ur�����H�n��e&�-%#2(�	 ��{�I;����@H��|QQ@7�d��.F�
D"]ϰ*B�3�Ş����ͭ+kiVo[e_��V2)�/����8�������,'��Q-VS�2�GD�=dS�8� �T�7�nTn�S��D�{e゘��@�8Y��%�k�M{/�G�8	���T��KxF���r������	�/e�����\�mM��"+������y"
�?�sڳ�95��i]�J���A+T��8�I�-���_��t�ӽ���ȁ��	�q��f�L�,�0���V���<Q��n~~t��Z1��"���S��h�|	O�+�y����B�T���h��!�K�ۆ���هn�5�bnϔ���F����\6ş�t����ڠ�����\7�V?�J+�-����J���8r��k�8#��~-Ѳ������O�����d��3bЊB�A�H�6kr�LO��$1��M3��!=3bA܃q�7ew��=)8|a~�=���ԭ�������(K�CR9熀0�+���BǨe���Jzj"a����{6o�8�VG�3�3�/�'L=�ɴ�Xsm<[��[���
r�)�8���d����W��kd���Kcn����Ou�2���]�1��x���U�R����ͤ��u��|��w�I^���y·����������ͼ�P�3KC�z����#`P�Hzv��"ʐQ�nf�\B t�&��*�o�Gx;f|w_�0�y�\&�$��}=����I��
�GN��a5� +Y����P��ᨪ��oeO�I�����S���ֈ�c��Y���@�����/�8Z�Ʈ̻��i�0�t�F��~���mka���q�Au,`N�U��e�,J�U�mCH6z*,��.�:X �=���i�C��k��чl��n͹��Dm�u�]LLY��U��近�H�+0k�O��ª%�p?( (R�~�A�^=���>H��:�' �L�G�݈����Kk�^��eژ�BW�R�*�n+�+�D\�^��]Ly���p�Q�\GF����Z<��,$K��B�E&A�^�?K�XDS���p_;ɕ���65�a�	��6z��:�a�\
#�_M�O����5������3�{�2��Քq�Nm)䶟���^L��O�Ć_�!-���h�UC��@dx�CuBռ
'���Ϋ������<�W�[%{2-D���PP���L�'��P�m��Y7?�}�~
����j������¥�������_eQϼf(q
�XS%%��my=hXi����*[6K�-}p�$8��O#[���g�ދ��.F�$|��J�(����"d�����$ �f��>B����	XTb�_�#�bQE>�f��.�$���Ľn�t�rR�b_I�h�O�裛�(m�ۂ�鶊�>z�e��6e&�3&e\�y�I�~ا-"&�4��o�:oF"��[�$]`˾HA�DM�) �4�I�uD�\
�|��µy=�%��ێ�d�R�|G`2��Yܸ����d�G��H;����*�,������u��S.��M�笾�
�x�wLW6cA�K	+�J��jHE4�d	�C�hG|�����B�>+�	��z!��r�g��Ԍ3�Yn&#p��ǋ�v�iX��`)~N�S*���3ʢ�y��I�ԯ=�`���g���B��"�Ꞣ!=���%�֠���eǟ���0���AX�G\�~L[����Nw�}wd�[�mt�^�N��įCK��@=1!㇀5�M�;Uq�ǝ�r��Mr_��w����w�CQ����L�d;�9�'��������I��B����Nob���V�}�
W0g�0��o�/+��GJ���1��T�B��%<�����	1E	p��.��@?��ڇ�����l��b
�+c7�p	�R�D�|d�T6�����Lo��#^���
�e��i���b?�5LJf~���y�������{�E���;^��PM�3��q���{"����mJ3iѢ��|�}�C�i	���d��MJ�����L~t�襋1�6L(�ZX�*�6 �^{������
�Y�H��8�����+�i1���[���r�e4�1�]��������A��y���O8m�^\�Ss�'���]�EC�Dw]]�s۝AYn�����/�扇�.�ȟ���������N��&�w��q	p����%�Q����I[cJ|θ?\-���˰�A�}sǿ�G"�7��h"6�h��9|��Nh;�}�Z�ͫ1�݊h?�C�Ck�YY�#�.�6��5#)Y�� �Z*{����Ө*s��+o�Ҩ#��8����f�z+a�q�-�������1���$Wc^�3i�k���իM�~�����%Z	t�b������kX�����ēލ�z��""5��m�S�l�q|�+O��ەf�=�1�e}�k�{�.ɜ��(��n���Ϟ��jCc��<��|:��{m�=���]h�����/ �U��ܷ1HdS_����<��5ڲ���A��g��)��MGt�"�/¸"��̃u�q�E�z\��Ϛ�(y���馩�<�hC��<�?���t7�\@k�-�Ź҃i}���)�"#x��s��k}�0ad�T�N��۹.���C'��/߭}>K+�'�u��X
5��(��:��Q�ɓc���|n�|*��q�2��{뵳��ح���b"����j�6��tT*��s����R
s �)�h�^�v��o
��c`���Ƚ�g�R9vRd�/�c�F/�(D�,�**�n9��l��n��ё'Tx�`�_q�O/p�R�F�vy��r�1��
��o��c��X��U=��=W��̎��a�|=�<�K� �Fn<�*���'�+怘�p�ӆxv��0��͋Q|r�e�x�؞_w�Oz|�}HF����c4Qʅ61�j��c���v�mj���_�F׀�^�s��УX�ŋ�H�".��
�W
���#�(A�|ް7�󤌙�hE�>�y����x ��<2�y�`/�S-io}_'f��5�Y��H��d�=�o�V+��]z/@�����)��8��C)�(�jJ�l��=��g�I��/�)�AtИ��j� 2ґ2_d���;��}L��K�Xp4����}�3ֈ?E�]�
�5��>���ׅ8�@\ņ�+��{JB���͗�;��O��z�P�ݒ�B�6	�� �7#���B��Z,8>]Ɓj1{�I��l?P���*W��,�ec�B�;-�,���tmq��	�&�N(ڹ��6n�'�d�'z��� {�w�|�����:؈~2��~p8�D��Rn��f��b����3�`6��H�i��3�)���S�5��r�~p�{�Z~ш������9�C!3_��2��SH[��Y����H	��g�{��$�m 0�)op	������6���W(Qτ <av�H<��$�5���l�(j�<T�&�k|����m�<`Ͷ�k�
ãw���(ljS�HOb�s��슿�^��V��l�he���T~Υ�Af� Wۧʲ�WŁ u+u)�]��t�H�G Z���l����9qsKp�Z��F��	��U!A�yg._�Fkw!�.Ny"���At�S�u�� �^�$^���hR���jZ�i�Q��J9[�~�Y=UQ,�}���D��_f;����Ʌ�X��w?O�_�v���mP�}�DU��&;օ�X؆�r������b���ԅn�'�r�p[?���OB+V��������`����h�.�a��w��n����mO?�1��>�U��y����,N��15����,��Hby�C	���Gba,�S&Y�e��4�6�uk�0��_�R�����#J���eX��J���9'���,:���A.�%ţVS	��~���cڳ��V�2��5���0hP����R1�QK�0�s����m���e�/��l �M4�e�9K2�Ѳ �?Y:�o��'����;GH�F�[��8mLq�.�3��t�KF�.�y��O��D�Z�|	TU_�r�[3�էk��_RG3Q���J�#E�_ݹ+cUa��8�{���z�.S]*���w�~	9�'��vO���6t��%-��@����E�!�4N��!'���#s?�ͯ�:=b�Gd�_��R0�
��醵Il%m֭W��sJ��)S8��,BX;��Q?e	��n$�Z�n_�9��Ua��4�����.mW�H�cƼ�'�&�@蠮K��-�{�[��	�w����uU�B,�����'���=\I_��r��7)' k�����2���� 9����1\-)X���W��6�<����S����IS��Pڮ�Ic���ER�4�H� �z��xr|�AI��!A7?rFEUh�4�ZU�_���V�`(�oIw�jӡ��t���of��W~1�IG�{d�k���z?�y{@��_�:S;�m�9�M�q��;�Ԅ�K�6�qP�~S�*<X���s�i�ZW��C�F��e). �~�|,�=��FpJ�
���da�?�3���i�̧e�Z���]��{����(��{C^#B���J�����	�<�_��}"�q��b��u�ҥlF��I�o'��q�{f��;�bfI %)�H�E�=�����v�x��+uv��m���`Y�C�#[ܶs��Ȣ���eJ�kB����S��q`o��j�l�\��M��C��[�q�Q���2��}3vj����q���a�ȶ��׳Z�_�k�����u%O�$�	s�[r'�QC0�J��[�ݥԷn�p���}z�,�4*s��(�*��ٰ��2��)�IԱj
�ٻ�Oo�-y���ʐ<{��+�+2P��Nэs`�"���C��!^5G9�.��Q3��!��n�OIz����� t5?ph�4�oDp7�j�x�v����[A�؟�U��Z9b�ރ�g��d���IF�[�M�-?�pڍ�MÀ�a>bJ'Wz�A�fB`_�BJ�y������O5��h��4ݎ���}�ݪ��D��כݩ]9�?�Z�@0��G��5��ۡ�dEO��h;�*<�ԛ!uUz�c̅��%v;�A|(վG�`�6��#,1�m�N,#YgJ^�.�׵�\Ll�TI���p�нw$�9����EV�ɤ3����W�u��[�\�f�a�o����Gظqx��xx�p���L}����������0��Z���<V3�՝�>E�������5Sl�����t�+�Ɨw�PцF,�V 7V�ql��onCo&�̰�o�p�2J��g�5	n`-1D�\����uD��:��뛱�*@$ޓ�c6���)�� \b�Q�9a(�;x���[GV�Y�����j���P+���tj
8��'G�]گL�.k/g2c�M���%�#w�
���V�G1�	�&�dF�&CgJΨ�%�w�.�lV��/���ǤF8��[�"LY�/�q֊g��kj�	��{k�88�/������v�tP-�KG��*�����>ȅf_&�FX�tu�zx���w	2L趩�PMe�LFN��/9/q�֙:�m���ú@ $B���8���r,���ȶ�Φ��R�~S �5:� F���Ӹǋ��w}0�$�:og���{^q��+S}�)\��!,r��`v��%����➘6/��3}���U2㐤�:�/��j���<���C �I��#{J4S�G&�~>�OJ��ǉ����>���	W��W��9ի��k�2�|6e���ݥ�U���
Jw8��q�@����z{������s)���jf�H^��HI�s����'����q��ui{C�_`���m�tʡ-�)�W
�"�C&� �F�FY�O���$��TV`\�Y�3G��>�D��Se���r��H����k���}m�+��C�~+��5ȓ��E�҄v��.�h�CSB��>��0�h����{{�K��,5��|��5�b�/��a��"VFu�B������a���w�~���ׄ��e���Ƃ��<u)��H;c�' k��ˎ �T�Ǟ���>����O�%�b��:�,�x��l���Qe*�&�������G��+rL�i�t3J�ة�/8�ޢ�A���Ɨ>L��P�C��~��"a�v�_�F��I����fȇ��<������!�P�xV�u��>\��Ouz� �C�Hd#V�E��uv"�3^�y}[\����wE?z��>\l���\����K��tt�{��*�>-�lA^`G��֓��H? U3C����S\T�y�፞���s�¨�Z�^#�G�-t	a���s,�G�S���