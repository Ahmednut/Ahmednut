XlxV64EB    735d    11e0�9�����٦و�{F�F�/u뻼��6��@j����p�����qP=T|ߝ��b�5J���4��-�-��/�r�Q�.�,�/6il	��u��|�J�;�X�f��"`�H �:ܯ�y����snd�I��ֿ�&;�� �9#\�͆[*5�>{�~k��[
.ʑİ��cN��Q��%j?G�j+F�b]���D���p�Ol��k�)~������_˥;�ZE7��%��0Sz���ϒ-����� ����Q��I�A)�g3l���'s�XȨ)BJ�,p���-{M�s���?0UZ���&Q"�Hz{��Qr(=F�&ڃF��f��h�E�a����r����9$M�rЉ W�s����
ᬅ;����v��0�B�n�I[z(�ksh*�G�ç�&���ɵ��NF�^+f{{:&��%u
^5��4�w��^"X�����今}7�R�+���\E�����Z#n��k�m|��(���"��ڊ*�ԄA�4��Xv(�4��=�N�e��p,��|�T���O�X�I�&��xƓ2� Q�;�0��ڕòXg^gT�OLF_\�GM�v�
���oC��淬��#��|�FpL�|{�6n��a��J/�U(��R�
��\�<I��E�A�����1��������8hY���<�|ŵ��+�kNK�x�~5�]��󜠛�5�-1J�:q�y't�.���*�T;'�j��5�a ���'qAT��:%I;R 
�$�߄��0�`8Es|��P��i�.ёZ;��Diٲ����|3j� ʃ((��*�VV];X���@6�"�`���9I1eL��-k��@�[S�|�n�Q���y��Cы<o�QZ�y��,0��x���WK�? <eB�E�j�9�Zd;�������JS�Q*��Д�%۬sX�0����٣HnK��i5�G_���
/�"��FE9c�ѧo8x���5(����c��!!�3���vd�~�VX�.��}0v#�����v�d璇���~T	|���G����!�e�!�>F��3����E�]:0��-~|��m��ݲr�"��U��8`�`жc�'�'&;���-�� Q��������t�Af<�G�7��{�o��.�|���Q�3e|��K~P�p��gx����Y�/�F�� �x ��� �F^W �i&��d$noV4^<W�D��w͘c�74f�(�(��X�u/����`G���z������K�m���?|�7����>�|p߃���9A�L<����}�7�q�|���1�4�O��%�\�%µ0П3�8�#��!1:<N�Yzq���c���.%��+�� m�e�)��.���W�?�=r]��,6I �%�#�n6��TQt;U�~���<�~�آ�>cY;�RҌ�����X{�|��/*'�'��ƑSE>�/O�a��N���ړ%��3WmW��u����U�Pr����2??��h#1��[�O�������I1Y��MS��'��?;�[���}��^���V�/F�$�j%j(�����B���H�Δ�幾���\����x;'����X|�F{��4�m�#��f��)���Fe�������i��co,���D��k&?%yo$�1�I���Öri�(`��{[� ��$�B��(�x ��cH�>e䴲D������5k�~־q��^�PA��aH�]c
k��jy���%��\�p�F�\9���*z8ł�����8-.?B6*w_9����%(�h���o��}4�w8y��ps��N����O�tQ�,0t��B8u�(�i�e�1�0��([��y"�l�iy{$3;ѵ@�to��_�GmrP��;����\��w��7&)��[\�I��C��]e�����HR�]�����P�cjp��S�=�0��@Eݎc{Iy�8��`]x8���k�ob0����MR������Ȯ��ky+�-���.�	�2-���`Ft�R�x��(f���=����8�+4w���8�f#������Y
��<+������n��1/OTa^��]�J�U;��x�i� S#�B�"!.�^c�)���0+�:j��so�J��M��>�*p�n�]q�i���l�)�?�&�H�E�_Ֆ�T8T�B���.�{>,�zR��h��S$k��J9�� ܷ
Ba՗m�)�����}|�hv���V���[��Q0��Ol
��@�t�RB쁧�Q�>f�a"~Фmw��t�i2����`k-��3l���Ln]e�"����;7����SR�zJ�ﾆI��Q{�"\D�kL�� ���*�����Np5�0��aCL���6d��%�e(�u��З%$fռ�(kM�c,y�����a�2�%�{1�������j�N"�)rf�tR
0�����И�*1���NR�U�*�!�:(��]��q~�Z��0gH}���槗�(EU�4'e*�h�F�$�3����8�匶�,WD4:R��zo�P�as�T'�7�[h"�إ_�L]���+�3��<R�����9S�6�f����B�2j�(�)�H� Bq6�l*�qd�B[L� �x��TfQ�!�d*R�w�9o����<*�b�
��W��=�|8��e��Z����7�A\�w�擿j��ڞct�3^;>��ҭ��-�z��l�o��)���M�\(3_|j���>��,M1��7�Wjw��1��ݮ��S@F:����k��`�	ԡ�l_��jS1�߆'"����F	Sժ�CK�� i��,��D̠���E�AW`��l��n4�'�����q^���ȕc�M:��=p>Ab�YN]��(�+mr�B��� ��(�P"u�ngwE]J�k?#���0@���b�@��|=��]�Fu��@�:L�!�h��N$QE̡�L�Z"�pZ�:ʓ��V�P��-�,���E�w����c�ꋄs��ӵm��� ���a�Q�V�%�-Kz��-��i]9�w�ƀ�>T�BA�1A��6�,��	�O�"�|��uE �GD��(9L$�,Qd6�P~�jL����rb7'�Du!�i�X�	���r���s:}S����`]_f��}����M Ա�^��#jӆ�a!�Նן��򃝃�	^��	}��=%�ϘV �+_��a����>5C"{|b�G
Wv��.S�(��I�pѮ)k��!�'�߸���k���Pݘ�qŧ��R�Z��jq���$L+�p"C��T�����#��ܙ�������w&��DP��M�$?�9G�6f^���������}/*H�����,!�g�VN,���2K9�-�� �y��o;��+t��X�mM5$���Zt�~��隖5�s����2;71�b�(�dԵ2j���4�������<ΔWm��p�8r��SB�e���4
ۓ�͚E���ޘM~5��Sn���;3N�d��V�#$�Z��?�|=��F��T=��3�ݝ<`W���_�	�byU�[��{uFmл��L�V�[�I���ZN����^@���l��F.��)ʼ��I��u���y�e9)W�z�Q��J�P��O�lWs+w�+��� ����)^1�̟��>�#d�"�d�_����eOȯ�=�B@pq��/�q����@�%)C�%��g�cm���X���藵��hf�[���Pf˸�T��#{W}��0�sy�O[)fPɷ��M��sח�<f�	Ϡn�����yї���j(Z)��	(��~E�]�pa���T�}g�d6���"�~�C�ԣ�[�Ax��.a��x׉i�e�r�eF@I4N_W�E����uJ�UI�g����e'5��c����B[䓅B��Ό�T���?�������\�	@��'��$��EQq{���5f��ʵze�,�[��)�z�� V��U6��[!�b�2���ܩ�Ll�)�ry=����	�4�8W.T,��/�⒄��x��
'��� ��IJg"�;Z�6��E,�� ���V���ʁL%��e�����@=�M�Ci�����V�n�9�.(A�[&����s��$;���g��M#@@��9g��$������( y��Ospr��&�]��lAa�[�8�5p�o	��:��١��'	��05&�r��	���_\�n-K�U�?>J�2�H��ڮ͂�ejܓ2��:�;�^m]��_�����C3�����8UbO�E�z8�v��~R���=�f��������-�w$���0��i�i葉l}�/����S�'�A]
�Yx���=R�u����-����b�5'"��e�$���>��V/��4s ���2C2� ɟ����S�����vJA�>��h�;+�Dr Cn�˥#����&���*�����l�������ix#^,8��p�&���ߩ����v�d?SH�K���Y�Q��A�{��.�U�i�7�:�` �S����Y{�*^�0X��d�c(����Pۮ���ؿ�f)Đ&̺̋�gH���
jV&�y//)�Ƃ��`��1Y��b�