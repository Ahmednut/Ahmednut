XlxV64EB    26e2     ba0$�ʖ���Z����>���O�Lu �)�L7K��x.2��*I�b�_._H,_h�cL��3{0�:d�7���Tu6ݸc��@L۽a	����3S���yDw_�[�~[k�[i~1�_T�K�/�-����0��5��pe���"�
�`�akR�g7w�*xS�s #+����C�up���]&�H�*:�;;K4s?�6SƷc���n�����I?�|�_����v�+DǬ/L��<����� �u\�GM_D�o�� ������6a�Ƕ��u)��qkM7J��G
)**s����3��x3�},r19�X:�ݼ1K�2�L�����H��Jt���4�1��� ��+�s���jJf�.@Z}J 2��d�5P��;�C.)��mg���ɷ�.pҊ:΢D�H�H^�:ۑ�6y���7�����tW����� �4�W����`R6���{����'�M�:c,~�����8�xw�Z���� �O\>G���2�*�I�d�R��	p��+@3UEd)���	�]~��\����$��pvEny��M@w��#�6h;�u��9֔=2ӊ���6~��G��!��8�쓄�z>X��O�V�4�"s~Weͨ����iD2j6ʟ��k4��-s��Xl����i4�u�C����y@D��pR�H��i�xq,$�~��zM���#�Pד�L�E��hξN]�)��/�_��^:{�"X�X�Dr���Bv높�r��-ۆ��91�,�2ɕ!Vbo�twy�!� y���/B���ğ��� ��q�xҥ
>_)��Ls�0T*N��3i�~�+7�	�$r�xb�����O  ��.��y����@n�[������3�<2�Ӡf�lj�QT�M��(}�=""�ޞj�D�W��#>C]�xr'�����9�a�B�{2�Π�b�8ݑA��lv�o�2VPJ1	�ԃ�P+��mޠ��Z�I���o0��j����{cZO��O����CMd��M�<��J/�nлА8�+�~�2AJ��4��M|����G��$6N;gÝ�-y!�*���+�/�H� /���]��m,�C�T�Ǵj����`AJ�O���8�:yṴ�٬�I[�2�7���LL��_�rvD[��rO��%���1D��`�&`bV��I�$��׾n�2�S�&h�[ԝoW��m�0��	�O���!��`�� �ZE�R����A���g�{�h3�'���ԣ�^'i��szn$w�7v�#O�l�]��.�[�����2S�9�>2W���%x��,�P��S����  �ʗ�ƛQ��$7_��] D�@�(8��N��t�5S�b3��D��[�,#Z�����˟\���$o��^��By ��/�}��$������]��3�t�M�5F�)�ה�t�-���$s���U/���$m�9�����Gaܛ��W�b�k�*�^��y�W~��[�B'�K�+F�����]��a���ouxX ����n��H�p��EAW�|���0En��O��r-��)P�-���oq��u�
�TVpC���E�|v;�W�;�4Mۮ��_41ќ?Z?�n
�hsg*��a�6�ذxi{<����B˲�I3���Jb_0�g�說`�
�����+Kqc!G�E:VwS��V��"c19���+�����BȺJ�)�^��B����xS�K,a�Qg�3���1���,�����Q�,=Aȟ��FߑM��O$��#��M�}7 Z��5�� ���P��@&�C�g���qG0x�w��f*�Պ�����lqC8%4��2 ���y\̫��D�F�`n�D�~}=old�R�}��fzNFo���Ż��UH%Lhz���c�l 5i�����R�F8t����p(����T�=Y�l����=�k �� ��e�~�e�;���k}�o�U��?��JJ1ҷ�%�d���	����ћ1�r4�U��WvSqu��Y�y0��~ל�E�M�����f�m`�)�+��ͱ�C"�`w�c���E������+_�=�žT{z`���AB�&RiG��&
��n<2��i�$HvBt��8�rW��@��57�l�eb�㴌F@Gδ֭����M!����X�/��O
��A�&�1�Y,�4���n��\���M�d[����'��!��|��E�����1)-�����RPzy&��=�����{z� �1&8�e��a�B���D��=��>:�X3�1`Z�v�H$��4��||�����m§�ǳ�(�^���L��Sy��3�j�@x ��rp�>���ň�࣊u%����A֎�g�W��ԅ����O@|�ȇ_�04���������L(�$ :�8���f�D �m��{�>q���&���G/�}ȩrqo��͎U�A���8�6�rV����[	1T
N/,3�6mkد�NI�z��)��!F,^@i	��5���^�A#u�]Κ����
�7�Ո����d��+ܴ��	5v�\�)��Jw��0�>yZ:(G���g^`p����[g^}Xv/ORFYѨ�R�^�Nq�k�Y�}��lG��|�x�4�HT�v�/N�TJr\FD+a�Y�����J^Z�u���{���*�s�zY`�!�TN?�w����_�h<��y�C"�M$��2����Y4�5G�q�2객��u��TXf�ѨF�H ��J��f(��=���*m���9[��D�z�C�
C��+Ҽ�������4]��-3W"Sz�	�6\��)j�^�-�굹AZY�������rgbD�j^�;��)�N(��K���
�fPgY�@�P��t\�x��$��ڪ'CR ]��:?�S��ܠ`"���۬��w�o�yQ_�]N�Bv��1�[�}M��ڨ6rE�`m���Tx|��?[�k�;�92�ܥ�(%���0��9Cr��$Isס	jo���J���5*��B@���1Pe;/�"��M%�^�