XlxV64EB    3361     ce0�T(X<ӣ���J@������,jttm�5�G�݉+��;;�nE���(�����0��������q~�i`�)̨��&��(r�ڷ������ʻr�S���	7s�C��5Qj�|����,E�2�������p|g��7ѣ�hH�l�K��>�� ,��3�Y�J�ip�<�t:*�zT����i�F�s�?<.D.��̻��K�\�Y9�Ȋm�\왘>�H�tbLN��r�]���`�JZG�I���I��;�AF��>�t�#%�<��HZt|Ko�V�?��B:U��!�੻96���͘v;�k���e^JD����7~����17�U���+�OӶ+x2�m'G�����1iDt���B��Ǵ���eU���#rh��T��'��받z���)ԐF�#{�-O�l�9~�]���`�>i:�X\ޕ���mD�DX�h�D�x��w�Lv��eCQhC����2�D����
�BYv�c���q%��K����͓��-�l4����M�t�po��S�#V,cn�OY�;ӁP-�h{c����WZ���9������?��NhjB���^���A�{<V���7�%-�U�����j}գ
{% �M�'�t���ͥ,,�
4;J���"�{c1�2�d�łF�'�K�T�Cg��v?߾{>TX�2(δ~K�w9�t�l�-Ϫ�)@���

Q���A�8ְ�Ŷ԰��G�g°IM��l@���B�?N�V����J�>cb
F��2������^�i酝�����6�PV���*�	��3����*�Wޙ4@��!Q��+=x��n�1۠�eu�ly �մ@p��J-��-�M��*���&1;��&�6�D،�Qj�%R��FY$$&�\OQ霣�g;�KP� �pݨ:zc8��_���c�ĭ�z`dY2��\d�wN��X��E��vn��^�����d;��5�<},�4}>l���-��6��HVƬ<�������qF˰S����Z��cH�Ҡ��_�n��T�K$�4͵/'���s������s��v�N�5��	��in{;��� <+پ��Xc�?��'9w��X�����.�9&�>��7Y����a��>Sh�������;^e��,��Ĭ%`��6�ُG��"g��s�� �~�u�ZH�V���.��z��l]X �bV�D���UgW�>�y����"A���b�S@�[R�d+@���Nkzo��qh���,�I�}� �4F��9����s��0�0iw�N�eˢ.���8+��8����]xn����*N� �_�K�b�\@�y���xP�`v����1;Q
�����4��8���~�(%9����,n�Ah}�Zw�>���������g��z��C�T�o��0OV�0�怤T�#\����O�h���F���6�8Bt:A$'2�+��+��<	o2�G^��9I{OxwxA/���;���j�~F��s�A�1E:��X R�GY�(��D{�e��}K�$�)����@|�[v�6C���"�[�*V�V���֣m�y��ԡ-���%�4�,a�9�fJ��M^L%e�{������>%��Jd���,s�:�V�$��Κ���f��a�,��XI{�2���1�hy;R�C�{oj�WqsI�����r�X3�N�-nb�~X��("8���@%�#Ѕ��)��X�IB��oʀC�7(L����� ��{����Uf�����0*��8<D_djK�_��� D6)t�Q��A::�fWƹ�B�M<%Ѷ�;���x/g�~5�ӰJ���)|��(+i��l%�tˌ�����J
q^#(K*��qܒ�@\mpN	ʞ�Gk_�����	��{ө�|k8�z���8ɸ�K�+�;&of�Y���4_�S�CeR��/uH��S�ٷ��"GS^M�6
F��3����c[
Z��+�3K-C!>K0tXMU=*�5������9,s�Jۂ��9R��5�%C(�V
8#�5�[-�������J���đ��US�E�cYW(�]���sbH�j�r|?� u�ւe�$?�����<p&i\/�-�;�<9�p��0����BZnXD��72�+���7�q�cd�e8�\LܷIZ(�<����\Y��{/��x���QGv���`s~�1_����M�&�g[�pf0��F&�^M�U�_���$����HR��C�}�n ���sM=�K����۵��$�rizG(C��v6z���~��u@����T����X��/,�i/�?��q.NuSEZA=�)[�A�L��ODJ?����e��M�(#�;W=7Bo�zڍ��,b�fo�+K�E��B^�?�g9�vB��&��ux���b��|'��(�����S�i�EJ��C"�-K��=����EZ7;�6�R�n��V3� �@��v6�c	�#�Pf4r��Y,����z&����!Ҁp�ID�u�g�x-�O�S4"� �8�S�0�����*Z�o&L�a�=�������'�u�g��Pc����G��*���etK�B.$b��֋5-��� Ҩ �C�v��@op�bW&�9N03�2�R��8�:J�7__【Y~����x۩���X���'l"��)���z1�T���%)���Q.kX �A,�o�; �K�v���[�C*k��FG5K.h%^���x3��"�w [ZΉ^T>Agv�:��F:�g�T��C-<@ârָ��K�ɝ�q؛V�WJ�I`,5ݡ-��#>}����,^�)Ə����R�l �]l�h�3�)��Z�����٭H��xl���D�R&XY �!�u+�9�m���W�`3�CU�2(Q"���/z�c�a�|鍺����S@��J��)o�X����)���f&�f�Ew��Ka���E��|L#�d���	��+�T�5P�NZ��Rjo�jM�j&��|z���c�����1�L>��<@�ev��B���h����y@-g�=Ԃ��%��H�߽�7�/1){$*�W����L�]vs�%w���$��T	���֒lgk��E�Vp�S��?�|�U~8>X��z&,����'��18UQzbI��8�l\��� �:�0��Ԥ�\L)���jQ���o_�-�v�w� �W����y�ܨق97��Z���\6&�����߾f��p��^�ipKL[=(eB�5�C?�X3t���.��!BL��,W⍼���<0N��ko"����JT�'h ��3�V2