XlxV64EB    1569     860K!+_�Y�	я;	��0L (�Ӎ��pV��9Q�����yL0��(~"���� ��쑂�,^׆��ڵ<�}bd�ρ��~�|�Ɂ7�PzE��5�d|�=&v5\j(z�� ���m68W,�t���hDH����nR`�����~r1��ޝ�`�'6�Mi��d�`�T��آ������Ŭm���uίҏq}�Z5����m�̽4EȦ�X�+�ʯU$(�&��+@�S���ڔ��69k�9�c"rhG�Ñ,�Scgx]�n��J���\yB�E����rG<)��;��Ē}�6�����J�ɪ-&�S������Q�y��P���Ͽ�\�T����֓��À��>��0��njX��rc��`M):��HU`�Cg�Mj>!JC!Lz�����M�<q��L{��5��I�d�w��`c���8������`T{�7�0s�;���r��1J l� ��r��x���zM��i:?8����i�*���g{+]ccc+�q��2�e��4����yӺP{jc��SP��<:;���4�!O����^��}�$�Y� ��n/ꌸ��±�m�3P�+���i+���I�vX#C�߲���YҸv��׆ȥa�����:�����u�E]�r��|9q��6���� :�:�!��ʻ%waJ�V�;��(Ð�H��V>a}Gyb(�#gB_�����L�|�9�]?�{֖���v��]��_}����-�1>&�{TM���P��˂ǰ�-���Ӓ!�M��4V�٬�Q�wF��̐��8�	�"�lDx'7i��R�we�2H�ag�E!�yo3�,�_�; �8Ai#�b-`��sxҙr&�@�"��J/.U�?6����������u��>��0��9Oi0�JiF;en����xb	�#즜j���lז�u\!c���
+z���x��UE���dG� ӓ���iɑ�q�\!͹���0*�w�a�H/��+�C�Yr�Iq�r4�SL{���(�b���������$���.�o���k�̹��o�mÀx����d?�6V�|�ߥL��`9U����U?�%"B����� 5�Jd�z�6��f����Gʺ�k����[�0�O�ފ�������$����N��b锑L��DT	X ��*,?+\�'<����y�Ł�=¸9�tǺl����u���"�?��4�X�d�+�F���];�r�K���RB���@D���G�|�d��wA?#�Y��^���R�;���"4�En($�)�ixK�V��3s�=ur�f��^�Yy��6Կm��?�%�&(DU�kz"��DWИ�
�s��f��7>634�#�s�I+A7���Fx���u��/ :z��T8*����aM|��+Eg�w��@�=0K�[�#�ǭ�:�cw����기�qy��f�c̲�b���ٶ�$u���e|����\Ǜ�W�*�+������&�R�%Ffhd�̑���:c:G�~<xw��o�=[A~�m{��E����	��@q�K�6D�h���<��k6>!�ۿ�mۈ-.�%Z�W�]py�
ґ����t#�r�d���\�U&�'j[���ڸO�|<�1�V�4cQ�Ю���9M6ى����Z8������3�)ѷ��̼��y�`8�"�1_h�g[�;;���m�{�R�Ӡ�R�	�2��;Z_�r�S<�%���T�,s1�V���N�Z��[(�K1=�j��k��d�=j�=i�_+��|fN�I,�������)7/���C������㐽��!õ\����𹍰
��O���#׽I�HJ˜�O���qH/��ϕ�6��7)��7� -���ێ5�������.�MNd���3J?V�+�&}�X�u�!��*�F�����\����i�ӻK����_I=0���+�Ȫ�갳I��r�z�Q|Y�.~��p�����d��m�{e��ظ䇐Q3���"��ݮe��.����wZ�6�|�S�b׺����dYn�!�\*�pA8�x�ʪ��i�gC3���2��&
���S�;bοN/���tӞl��N��L�
Q��?�*p��5q+D5^
��ܚ���"��/���