XlxV64EB    181b     980�+~E�@��l�B�bt �E��] e�c#�Z�}������	��NH=�9�
���x%#���F!��sWc��U�LmL�8��_n�l�g���uC�'
�_��gd�����G��cY�M!x���!��Jy�F�pM�;v���
i�>�VL����2�HkBE3ؿ�@bMϧ�@#|a�#�?� C]vs����o����՛�.+m�X���~1�Ӭ��l�������Wb�E%�^���	1��ob^��|�
������@8�0H瞢�#|"���َHy(jnNp*������-���|�(f�	ꄗ�� S�9E���<j����ô�S���W�'7�T p�ڂ�	�8�	�m�2\_��(�A�	>�]��BP{{��N��G|��=�����
��Y^�1�1=�x�I6i�C7���ljGֳ_��0�s�b���ڷ���w�Uf��b㝡)��
;*!1!Ƨg� �-S��~�o�^������.�e���-��"�J�T�''e\�~ݘB<ȇ���>�J�S�q.�����\�U,j��
��;��٤2�����g���&i�)3\S�]A�X��0��&��8w(�0����F�I�d���e0�>R��6iG�<^-���Nc��y�g��I�D+sG�,�ߎA<k�THqe;0i[4�ö!q�ΰ��dڲZ[�nlV��Br��q�j����ڠ3�a�i}x�ߞ�D���fO&�{�����xa=P2ҙj%&�;�#Č��Y��R��l�6�tH?�	AX�����>�,Pj*�*���� H��Kg�(�B�����q�%� �n�en]���\�����$����\~�MY؏�oK�NvL�fO�`�!�0D͝����Ĵ�H���D��eQ�A�a^��|��V-�����G���v~�<���{Ue�h�B:��L'5���jG�� �����v"
 �LxE�R�qX��d?&|6� :�+���~h����[\��k�Q�#x ͢�ɵ������N(�\C�y�8�l�Z8ݛ�
�;�i� ��&���'���Ҁ��E�0�p_��UWp��_tA�~2P�������&-^�޾i��6�������Q����m�܋��a���=P�~������5v�xZ�{��ܺg�K���W3�z��ξ��Nq��@�}C����pC�������{--���@<; a,�%��f��\ 3FP/⣍�gؒI�Z�t{.N�Ρ����RQ��F�EG�qR��T�HEa[�hJ�+a�+��$~S�����Z�_�N:`�#��\�sz���ՠ}��c�����C/�`���]�.\U!�X�/�o kU-2�����X�6�xWFڡ
aiA�w+�BU�OK�j��LT��o&�z �˥�R�yD\����d3JԚ'��S~�ȸ�4_K�O�d�k8��Û��6���F}�m��^!'.����5
6����������
8��*"�M�
i�S;$�dT��a��*:�f[Yt_��`p��Þs�Z��0���6Y�{]q��
~����G�n�w���7�41D�u�?�L֟#+L�7�a�%�Q�</�8��5p�e<x��&F���V���cR E5�����ch񣲾�}a���gӁHӹ��P��Ju�5M>��8� ��F�G���	z��	����R���R� �LQ��,�wM}SE� ����v���`��o���K�ѕ����l������gA���}Rkۉ; N."��/�IQ�c�mq��j�H.ϧG��U�f|���2u�TWl�K�����.������%L���h��2�����)v��+�G6�e�	�u%�S@��OQT������b��(��f�*�p)A%-�xS8��ӳ�p8ꢨ�` P&_�������`I���")盃�����"�ղ�|�_ha���hQ����Q�㳽z�G\9���S�r�&{`Q)�ybڈ�Ss�ξ�dZ6~K;�Fs�eSvK�`�z�٫)��p�F-�)��ʦ>zV���-�s�f�r*��Xu��1Ri���E�E�@�9�)܁��������V�����?�e6h����.���fd����X�v��x D钒�a�}�Y*A���aW\zkjq���i��e"Q)J��ޥ�J<���|w��G��̫�l`*x.�nk�2n��:(<
~�`�bw_KR�÷�C'�������t�G3��N�	ΎX�H+WC���g�k�W�W��O1����1��U'��[Vm����5^r��T�v�Ų¤�o���]WpR�O0}A"�c����xc@t�a:?<�2r�L�X���mx�7���cI��i��v�('I�(���yF�