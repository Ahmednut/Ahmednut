XlxV64EB    40cd    1120���.Ѡ�+��C[��Ȼ�ڄ���m���!���r��*���b�ٟD���M(..��V�b9�?l�;{a��B� ��t�����`��2�����*���d���6�����t{��������0;Kb��I�
aD��>iEf���?���=~�<R��b�6��<��h�֘�[W��Sz���⎐�1"����"*�ZZ��kHTW���M�æk�h&#������вM�r�$��n�*bZQأ�S��E�Nx�w�گ��=p���;q���[�*��D�Gzҕ7{�ޮ���Dx��F�P*Ѿ)���%s����i�*�`�`���C�9$g;>��pa0 5��z+���Y�ȇa��ʘڎ�Q��5l"�]�x�I6Wf�mȱ>TE<���k�4P˺����:s(�d,!�A��2�_����$-���z�Ot���pp��l�g5`���pcs�l\`���r��\��<���w���Yr��=W� S��"�5�L�<�q���}I(U�]����ɤr��}�n7k���H���Q�F�զH,���T���c��0g�j:v�a,|������m��- )��GM�w1vr�k�	��~�e4��G
�eowH�S5�ª��e�Ȣ#Hb֫�X�`Ɏ/&��tRK	�I�9���m��O��c�~,�i$���y�/(�̓vH%�k3���tވ������/��p�J��~��;�Ěf�}�Ҩ��ˮ�"�����n�}c�!�9��~�Q�­����m��L i�i�[�q�'���%[�����_�6DB�^�����S[8g�-t+�5m�\����Y��P�@/�"\��G%AR��v�F+RG��=��5��f9ؖ4�jB�J9?ư;[X�!%|���]�]�2)��sƂ�8)T@*�R�)C���Ě�@�kk��m+O0ُ�Pdz��Bj�D1+���)�r���Qз8�����u�-7��������ª{RC�U�2�_68���������.x��o8xL�JeHӹf	&�&�b���c�Q��'W���ߝ�RyS�5�z��G�=1Lɯ��?��X1�����'ާ��k�L��|Q#կ�!h����Q�V�F"#��eM�
�n7G�B���)y�ڨM�\��|x������
�ʕ�����ݛ��v�����R��VF�If�2ҿ?0$Ͻ��EX2��fy���L�|��~��I�����|���aTכG70Y��+89�_ԍ���?w��:8`_3�D�/�-�V �`q��!�U]��@�Ñ�s�Z���@�H`2:�x'QhϮ�4��}bK�b2Z�۠S���K�D��!��ᡓ���YV���,Ii�20���*~�� n�g�o�#�f�Η �z��BLI(|�Bb�Q��AY�O�9�7��.�3E�7;p�>�G��9�P3t��FYٱ��<Q�v�o}?0B	���.�<�1Cdbh}U�?���!�$|�5R�KJ��"����� )A����a�/-��p/����p������zOu*4��d!��v��A�"˓�:�Ϯ�
�m3��F3�ch�{j\���e�VW��I�"��Zx�{n|�}�iy���Y�_\aM�X�0l�J�(�J�a��f;\u��o�5X�Sp�����}��'L��.�[��9*��Ȩh�����-�.��\����U��B=��jr���ݬ��.tcaQ0cx�	)�'��e.Ԝ5Ƨ�ONu!���'�x��R���bw\�Gƴ�׾|ƭ�]ba~��"�Mz>��l��#�2�@g���S�>طp�;�\g�켥�����Z���$�J�u�d�,��rO��Ч@T��k���u��p�'͎k�*�:���8����E��$��T�fͲ�7�Q<��B��]���;���ȱ<�
j鑳���/�ɓ��[�)�G���۳�pq��c^�<|sS�M��$�r�F@3{F��Q7�#� ��x� ayZi���rh���y]N;Xl�T
:�(��^�j�7���P���}av�]�C���+�W���ZLX�kZ�����G��E[�w�׳+��q��'d"f玽
ӏA98)�k��A3��8�u�p��0R�%B��y��H���r��G\afr�W!�N+��w�=��o����Û<C��z`p+�p�`A��+F(l~ h����d)p�B�9z��f<8spN0�[�r�N�濴�����TrM�f�C��>�vΨ����E8����R樮�Sw�+Hw$��`�d�&�~��,�LB��������W�X89�������{"+[:�JQ�Ηxϓ�sTL,�^��;n'䊎"��Oo&o@��g���_�#��y.�,<��\e�B��
� !j�Z!��f���͑
rq�pU���!x�Q?C�?����&�D�w���t�B����k $J@��'�k��tFr�>ѱL�b�Z�vlW� bK���[aM�]L�{L�D	��3���Cg�乽�Z��fb/�ձ���%!:�\��+�j8�@�B0�pe�X�U���>Q�I��h{�
H���7�q�ʍ���)�U�j�*؆�sM���i=�I����[��dm,�_	q��e&W�V���������.��U���z7k	
8�6S;���.
*V ����]��W�n�B/Q�:2��I(k5��m>6Z&���:>ܵy�Xw�
����˪��˗a��ڷY9�Ќ��*����&�� �P�d���ͪ4=�K�y�21���}�z�˄��	���'�=..���#�m�s;^~��֡����^ ���p7��G�40�ts6�t[_h�|�%~%�6�7@�y�w���{d�Ny5����y��Cj=R23l�����Ba�����ଔO1pUV��]TD	2����m��+�
�Tv���1/
�����7�(;�,v�*�'mĚ�{�[֑����^:���Bϼ;���x9�� �K~�?�}/G�%�%�f-�-�V�#���u����5m4�d��y��[�vǰ���_\�jiZ��?=���al��c��=��w��6] �^��A�0I��*��I4��,p~X<��Ӳ��KR�K;�K;AI�j�ՃQ�Q�'�0���1䩆q'I7�S�(���������o�=����W!~�{�wI��)��� �j>?��y�jƱ������j���a�r��Jz}͖�*_vE���Ժ]�ij��ҷ#����ׅF|o%J��~�����?4�PD�P����ʎ=n���g��)�p�*	�^R�J���L��9-�`�����h�&i��D��ră�X�Tn��	�;�V�v�]��)_�;��F�d)5[����we���$z�r���NE�m9A��PX0(�}w��+��W���.�aT����� q�9��t� z��O{I�+H����	�ӏ.�&��w��N_�F��_g n���`ع�l���6͏+��⹿�1�w�-�=����L�)�j�I]U�8������'6)��lV�^L�L�������Zτ1#�TV��@~{JӮٯ���[�3��%W���g�������A����T����.����6�Q���/��"��ע�<��#=���.�S<��,�	��D�c��#w�pI��#s���t8�[��ڝTgC	̔�:ݿ򂎵m��46���(�g萼H�E�e=P�}ʽ�hk_�}|���
�`����κ2�rq�9�#�`7�QIIX �V��������g��K���;n/�I��)�H�������BV���!9#�Ɣ4.����[~�LxׂBp����ְ\V���Ht��`O��o��\FU�r�zl�a`ޯB���Ѐ?9P9�9+�dA:��37���R�]����A���ν�t"������KMȊ(g��
�&�L���y��ܸ��O��y�r��L�|�~�w�뚳sPީ�I���C�������l+u�P:Âg��% ܺ����^�$�3m��
��p%�����Wy��>4
ܑ�y���N��'lΟ�f7��Im�膭��)l��2ve;L�6��jˆ���۶�_��W�����\TB!�����`����J]��	�Z'��<��f�����.J���2HI\�y�l��^�%=����N҅�w�m��x�2��Gh��'Z.1j�eR`��5K��L��qr��/EDB�v��ϋ�EQ�"|.C�5}̺�h.t�[�9�Ų�Hf]�$��Y&n�@�f�B;06z�$(�C
cԄ�X�NqjW]����F�O��5