XlxV64EB    fa00    2f80���* ��ɽ�_m�NtDt�]_�SOΓ-����g��0~U�̠Q������Z�h��a��(J��){Y����q���S�����vs���H��B�+{."m!���_�x��q}gv�!�J�����r����T[��(�_��x����T. �C�s?�����C�+�� 5��`�����bc|������I�I�[�����z���<�N�p�|,3]k�k=�ٛdm:���Ie���T��Qc�z�;/�G]�����H@p�q��;n[?�	5;�6 Ӌ;����I����[�yb=�'/���r���r��x��'�P���(3�='T�n���N��;O]��a���_\��d���_y����+�g���'}
\�>�э�_z�sOh�L}e�����u{h�N���X�e�q\u(�7gHF<��A�xF��Y���9k6���55ÎPw���`��D���	��
P/�����k�[2(�2k8kE`{v�Z>��a��^8�č7u?9�z\v������B^��aPO��(��:�KߌA�J8��`߲�Ҭ}��Yk(
�{�����>z�V ��na�EI�وȕ�����2�?�����%��,`�w�c_,�j��| c���:~�mk武�ӍI8�h�����j����Ak-A 7]~��Ș� {N�՟��*�BM`���lk��a�Z��Id?ӷ���uv�4tE���AT�5��M��씔x����%�`����.�k�%! y��l�������S  ����K��S�J�	=�^\��21&������� ��6��}�xW���� �T�7K��{S��m`륱�'�rn�}${���FO���N}�Kc�X
`�T��U���3[�]z��b�j<�D��xo��)��g�B�Ӊ���-+��J(1�4|�LR3Ǩ-�u�C	f��p�̍��O���<59���+i��}�|�a��m�z�B�k��=���=���#)�>�i�k���&������^��{�9J�7Q��8!�Aӳeobv���G�\�e<�vV/����R���oi�o���ْG�1d$D��M0�"�]x�Y�vR	�+��[Ƽ�W��j��;ße��B�.�eJ�z9��w�]�7���/�� q�0yL1�m�I����m�v0��T \��,��U���
�O6^Q^��<�D��
��4Hk����V�|���_~��YD�����]Cy��\FX�?���V{v)����/��)��5��Zۖ���VP�O8�C�ZY=���p�J�T�T�9�ʵ��9>�����f<���e���s��T$W<F�~P�(^x�����=&1	J�rwx�-��,`Pďӑ)�.�=�(�'�sT��,�Z��e!"�����`�B���V�E�Yو$�c�q�~�����@8ߠ���t�8�t��<�U��T�_��j�/!?#�%���tv��cTK��xC&4$���-
5���x>r9A�H:D��ٗ%0ǱS�I?���_�4N��4�a2w�Z!G�5��Κ�~�f�C!>�X�㵁�ݮ�����f�-%��������\U�C�U�D#x�~����߽#�!7�԰/=�K��.ĔYz����L�)�-τGܴn�#%�F¶Y����Pv��aHJ��p��r�:t�C��"����8�{߇|���4ڪ������n�@0�/��dܩ�d�{���F������R5/���uR͌ԕ}p�\mSU����Ls��RJXAx��K*�L5�'���$[6	�����C�� �I!.�#ЕR凖��~>Rml�����-+Nm)I����E�����1dO�ڧ^����P8��AF�@�v�O�$��.Di����{:��Yd
mc���'�49l���y\�N��c(�u0�?��jt�GN�Z��|w�Xa��=#^d�fOCQ#�U�4���į,Sŋ8�ѳ��T�0�r؀�ld���a�����Z�΂��z�9�}k]GL9`|Y�c�Q�����`��w�6#bj��#� �ەՄ~���d�X�om{3}���b��p����F��Fʣ�)��0�3��ʝ_;�5��?V�����r�!��.t�Y���9��$M��y���}(���5T�1I$���kR�O�ε��(�xqU[���a�v寨����Ģ�D �+�{uy��/{�Dj��'��gs.��S�2�uw��K�ȩO��gN����NP�1�^f��]q�<wl-^�������
X��<�6� ��*�!�Oy Ϟg�+�!���A�To��`�R�t� ׼>a{6p�Ue��*o��6C�B���:0Y5�W��_�����'�IH+������9i!
6}�Jr�8(phͳ��.c�B̒j�O�P���ia-�� ��
~�IH��㵃��N�
�RQ��DR��7������q�Z%���'WJ�2���,z[�����Qvܮ|'+�W"T��{� �	�3���6��63v8�s�E�&]X�03�g��� b���-x�&���d���3���J�s�a��/��)�F��B9D� ��U1���Q7o�L��w�,����^����q'כ��2�ۙ�[���'�����Bbzm�ऒ�a�/'&e���ڛD��a��(�@5wɽ�X9�X�h+Q�0�kL�����ń?q�1���t�Й8,���aˇ9؜��A�L�V&:��13GtyU6�b�hb5�I�Y�c��n�,�u�cT�!�*M��cRy	�e�?�SJWn��]��ty<p��k�,48��,\< �;8Q4��V4D�7�Y��ݽL5��x:��aB�4��Ŭ�1�}���������(�@O���<�l�b���*�� 3�^���N3S@F��1	-�u���7甚����]}g�M}1{~>�dU��@m�hQ����<�����2��`뒗���O'hwNե#�GU����Y����C����l�L�b
ӈ|���t�	�[�,���� #���fXZ0Ł
$��	�m�p3N�T؊�
��V=ȓ}Sz���ª|{F\8�'��Qm����$�1��-]���e�ii��,�8�@�n2�V5����!I�m6�Wr�Ȅ�s�H��d��k�y�'S��@{����sJhF�}�`�+(s�U1g�g�4#U�Ho �[����n���/-�3�)C��ڷLk%��m�e8w�Lء��s�Ï�J�!䒔mϵoa����8�J��7$�}evw2��{�{�PrpN�z[`B���Ll��=�'5!�`\Tk[� �0B���]
E`�op�0G �����ԝ:)(mK��NnI/89�t��̩u��0�=}�?�������Y��ji��}�Jșǀ����">/�*���p����cr ��@f��k#�i�9h��P2�|1��bv���fT4��A����g&m��L�|_�H�O3�ܧ}����k=Ľ�_K�z�Ke�3�+�1��2� ����)Ss6�� ����%fdP��j��n���H�q��)�,ZX�3B�ٹ[dy�kY�$�A~��5|#z`��F���c(0��"N����2R7�Jэ�B���_�0���YbK^��!�\|��b�r�I�|��?N�eI=H�<r�,O�j�Ô�gAbʡ(C���s�v�\���G<��`2eB��SZ�U�La���tqj�@��s�#�9M1�SwS�
/���Hb
ŕ��ӱpKA`�kk$w�Z�XXn8���\ʱ����վ
KT8c^y@K~#�>,�.)g�/��*K���d��se��i��_�/���c���Մ]3.��Z&��ezi���s,��?.�=�����#�����3�NO�=�� q'6�.�<ޓr�)��j쁐I�+tغ�k��kJ��R��h�)L�N����%�b1k�17�*}}��k��-[�7��\b��9=I^M��qs��&|�7v�+�6�]�!]�r5�G��[���g����p��{��ّ�ٵ�+B����</曵���6y���j�dS7�����9 �3��im�ߍ�, �����O�A�Ky�'('�/�~%�����c��b,�0�c�D��pݐFC�� 1X�8�1�f�!n�)���_���[��P��d���e�&�)+8��a��|������bN�UF����Kԏ���{'b-��VXk�`j��|��2�	����mf0�v&�S-�(u��!v(��x�l��r)�Ftd<b-u��}#�4��.���/�L�����C�cl�t#e����]+1��Nzk��}�}MY"�}W�`�n�� 4<�H-�����/� �����_$`����� �c�*�P��� W(�v�^�*�+ae��j]-�7.`m�aN
����uę��C�����
]h��3mAw����U������f��{a����T��r�,c���"R�c!�.�]�V�[<`�C�w�<�DG�`i̴�7�c��.��Y#���\�N�4`�j��	�N���/T����Uj@�=�*�x�)�Jo;�f(ѱJ����?3�-�+^b#�OЪ��NU#��/�{�S�@9�Lw����,%4� z��OT��vF��T�2��?0/�@47���i��'j'�È���шϡ����%D�RM4��P�H��:�����&�>:j�습'm�;ޮ�]������&�
�_kH ����أi�h?��S��C�t�D��Z�)e��e�%�}��;�,aژ��4?b�����6j9�6a7ƴ�397'����e���8Ͳ!��t�~�"�ۗ�|�vlJ K�-G5[�MD������I��{�EݜW���V�w�q���6A����A�8V�P�4FY��B��#�H��#�����[������$K�D��o$=x�Ґħ1x�4������2&�S�)JxTF����t�Z�溊j��4�=3�~�}C�=��-q���E���R�{��H
��Y;S�#(���*�o3n�1�Kn�q�8���V����ŋ��+����림peۇ㰊.�׎������!�����dm�>�>���*=i%.
 ^��Wlob=|<_����]���O/���[NRr�W� �0) �)̌�
����,S��"�d����)G�f
L0�0jq�
�g>uBg���܍�M���2�ᚐ����R��z�G}���v�O0�@�����~��37�	�˾|͞L]VLp&�:d���R�D��k��?�t�0&+;o����<*T5�X��l<(J�ԼT
��Zm�`}cSt��"�ս  %B�.��^P}B�	�G-�˰�X�*3�w"�ٓ���$b�&��DQ)8[[AU8F���d(��L^�Im+j�uE��ɫ�Ȃa2O1�Ŷ�=�DJ��]���A�~{%&���f����U3f���+�B���P�BEd�98���9E�,F=�z�[@=�H��/�ﯢL*Qi��j��NK=7.�I�b��}�'b�D%��!%�7y�q���t�>`�۶6�U�@�y����=�(���f~N�I	ۅ�<[&����Fo/��7U���z����[!�%������^p���J��י��"�K�����������>i�B���'2��_��IS->OL���2e�(���Yw�`�ݣj^��>��x��͆�!1�h �B�A~���8.�ˡC@%�����կ��)zU�r,&o2f���Jm�~4�%��[1hp)�h׹�#�����Wy����H�or~_:�l��8���8���hGb.ۖ�7�x9;]JZ���ha��������S*N�`Rdg����X`�.>�<�h	�VQ-.� �c �?kE�Qr��1/�T�*g@|�(�L���C�pT�;�{c��#xk�!h��.�RIB�������K��>Z�:M)U�q��c�aU/w���T�ni�����%j�h�Z��Vx?W�^���˹���/{l�~�Q
�?�J 6P3N�Mu�]?�=�_D���5�=��=�v�ޙ�h��sδ�X��,��M��c�8~�c�`�v�q�F�kX�<�Q�EK�^2K�9�4YS����Q��,l��wE�X;>~���@;1��o1�'���-�..�1m��cA��<,���f#�Ĕ;L�5~_�.؛l�(����$e70"��<!�c,;�K����ț���9�z��[�����^�S��t75����y���J�w�%�L��_�n�d�����]��7��K�t=���j����N8���{�r�^��8Hqx�~��{M���f�Y�^�����i��.E$B�f#C�)�c�"��&�
x��Բ�}w#^�<����3k8`�����m�
�Ы3lĦZEX�r~�vq�ǐq��W�c?���_َ8�n�9���V�1�j�gɀe�m�5E'�r�i��2X0�.�v�]�<����]a��D,Z[`����Vcl�����<����jD����U�G���R8�pp0�S���gjs��X 
�b��M��u��~:uA��`PӟU���;�Ӂ|��oa�&�.i(7u�4d�b��m
�-�Jd�g����^!��"�N~��ǵ�^�7�+c ����[��{y������jF'}xNg��'h�KM�c���N�BZ�1�4u4r�kX=�jj��YüC�td�
�XVg���(κ������ ��=�@q�j�kӾ����P� ��Y8H��l�5>����Fd�U+d��n�徲���F��Hiq���t��AE��� �0�h� �Q�H��cV��A;���`C����Р(�������~hh��"���\{2i�
�d1�����(	�	���:���*m���99�����5�q֢��'����E�c��;� �ʇ�Z��q�n�x�/H�Wuu�28�\�Y�U� ��_/R,����W6KAt�-F���3T��_��&�TYn4*���$�S��f�͝����X5Ӫ=��nY����Ϛ����4(��ӌ��Z�ʒ)]Y;W���Iǌ��T�D]��xy{�]�� ��ˋ���W>��s�����<V�(y�s��g�����p�G3��z���ٶ�,j�6�Yd���xFU���^P���7�g�b4A���u�Ƴm�%������o92�&���� �@��Pd���j���W$V�EK-�k�������ڝ�]s!��d�SFΆ�/����6��8ѺX�'5��M���`���J��t�XY��#���L�O ���=!R�eU�#%�C���M���c%P���2!��A������J�� ��cjH���vt�HV�Ud��B�G9���Ά �s�I�	�i��J*z!7�5����sh�!)|qK��ӵq昽
~���H���Z�E�9P�is���>��@$��d����Sш�C��>�;���� ���u�5V�\e*w�����~�L=��EL߁�}��S����%y��+	�T�-�1e������C�"E��h�u��5A���T�gM0�G�<����70�b��(��b�1�5� j�cU�M�;מ�f�� G���2�5��� �X')1?7�_��o�j�<R�ro�=���V����%w�T]U`YW����hĵZ���o%�1
�8�γ/,1Js��N/�o����{������X�ˍ�5�t�p������)w�_��d����c��2bQZy�Å�L����F������f:tDOC��Y��F�n�0��^�j�yI-NQ�����ɀ�������:% e �m��Ls���v���矣��d��3S����F�^0:������1�+�@H���٪���2�O�4CZ�4*w�����&m��H�t7�Z��k�ԡ,�A��-�7^"��o����@��l��~�?Jk�z`�����\R%�	<�`mq��I���zcq��G��m�w�
��ቸ�ˑ�+Q�8b���h�]®�`�/Cc5�L`�+%.%����,Ո���D�'��!)� Z�����@0�־����Q�5���g�߸u�BϿ�p2	l�ɖm9�Ԯ��ɐ�x|r�%x��2�K����$p�z�+�?�I��[�x�Z�0�$+=�ɉ�Ӛ��ư���O�hJSd'�45i�|�&Yߓ�����k3�̂�Г�%� c͙�W�{�)N�:٢_K-G@ ���"7b�,5�����B[�b@R#���м	�I��R5��}��V����˖6xǓHi+\$(j)94)�_�y���ЉPJ�������V��,#W�Y˘ْ�{u���3��i55���-U%R
��!ɐR_�[�iҝB~�n[�탣� �D�ΕpӣDv]��+�fg[�7�;��q�8G`u��{��D�R��]�X�P���&�,��d�F���	V�*zW����;T�X��>�ui�{vUaǻ�vlI�2gD�ð�L{(eH{l�����ɣ���#��"�M��\���+{�<U1gʱ�4�rW}����S�]��z�!�T0�1���P�N��/#L)�,<��>�������]�|�Z��݅��6�������b�բ�.��C�^���9'Y���T6Jc�w���uĈޔwjN�jH2���o��-_�#�F��f�`sÿe3+��#����O���+��������d�1�^����*��'Yo�9D�k(M�Rsx����"	�΅�_8N` |�͘��,ʞ^��r;ݕ�U��+�lC����v	
�URj�V�::�ᮿ_MF�rl57O��9'68���pA�^V=��7o�Py�Q}e���Q����	��{��,�C�۱ߞj��dɴ���oꓟw��X�LK����e��<������$d����	k�sZ��O4|�mFuW�۶.+���i�E����!r
"N:!|E���l�5&��@�Ɯ�>L]�թF�lΚ����7�&�`Ͷ
��a��r�$���:e���6/�o_�*v��~B�ȩ��w��gȰ��8d����v� �;�/|ì����i��ʑ{'��h��#a ��ʂ���y�cY�"<�b>�O���/nVu���pH��ܩ�%0�ݕ���Ёj>��hP�>�Dy��(��Wa�$9��%��1$�^����Q�typ����D=1����'�欹IQ� o�~,�����O`E���r�H�|q@��gxL䊍�4Û�;1FNFq��h���Xe!���=?d����M����ct3,����˩^���+�1̕~/6�X��F�C5f{;�3���	�T�o�V�~���N��M_WW�������V4Mf�h����J+ ���ߣ́h���9������L�^Sbi�r8��j��#��B�~r�p����9@/�c���`��a����e�T�����I�q�������7�r��aAtW������P;���ު��������8n�Z]���W�Բ��~#��JWA �:<�(��?�uߐ�p���PvE�r����o��{Q9d�2OSÉx~i�M����d����p]{+ek���i�@&'A��Gl�1�n�I�1�z������ӻhȏ<$��h�����y<��9-���M:��5�� k[Řo̗y����H�洱�;� X�
��aP���W���y�Q�Û������(���>��7�*�(�O�f�>=ڎ���&�#I�؆�]#b�����Q��T�(��j�g��x�kI'8J;����-��~��Y��������+��y�w��r~3ĜV�ᮦ<h&����%��(���e�V��۾�Ĭ�.�O?��z%I�B�P�M�������rQ��?F���S�������1�l�f�UT�[;~�{��X��6��H]Զ�y'�E6�-,%���\�Ͻb�r<�ȃ֤�����D&b�?�z4=�Tܩ.���v<��(��%>펁۹�0��Y}�ؑ)>��I��I1��ҋ]�Wo_VX8p���R�'��F�A��O�=J�ǁN8��k �qI�֋����h��&]ߏm�B�$�V]�'�Ҋ��0�a<J��uD����mb�����[�8�7Ը���)�v��1��l��]�� ٩_iok�iK��7~��Ԛ�y��>��I�o�� 3�l읁lS@N� ��[OV|�9S��\u�	�9�6��K�׳��2�B/`.��}�XN \G�Q�"eڶD�ec�92��̯�xn���S,5w皔���'6Ң�e�������=y8U%�JP�=�?3�ZT���qtxK�d�zc�mn��y9o��˗��/�����3�Z F� �y#1�r��V˯��n��Sӝ=3���~�b\^Y�S��!.Z�!j���+u�++[	g#�I�ޘ�����58���K�z��E�pN/P�P�e���Q����d�{���� �*i��Kȱ{�3 �P�}�԰�
຿&��o�KiSѩx��V��l�&3"Y�/��-3�ێ/^%�N�����:P�<Q�!�R����m����*¥�K%����)#ftI�[�i�1�b��V�#U�����E�k�g�����>� �W�=��êO!�ƃMHgjz���ǛI����s�� �����Z������[���f�S��9*�Z;���8p���7�*��OР��G%. ��v-�j���q<��{K[�g�m]�I�8��W�J�ѥ�^gT$����e�i��&@,�K&���P�{9x��5�)���(�!�f�Bm��k��5���G�[V��/�MT��h����[~x`nyHR�+|ԋ=x�`Cy^�?��༡�|AxU[$x5��Su[6��+ �d<��GP7�qF�8��G��;������
�ۋ<�R�"ϮI_�C>B1�
�w�8^�=�ng���<����>&f}~<�R�\F���(����#���z{-���kFR]I8Ж��x.���pT�)�n Ol�����;V�&��M���j�WΌ>�1�Ѯh�8�Ϗ�YzG�� 1�n��ιb��{���`zb�S��ؓ��vA��h��.^������+�o����j�;tc��^nǨ4�0Хx�;LLbQ\���L��R��C�@o�w��\5� �����t����@�U8��W�

$T ������c���i�[������"D��o=�c�~ia��jX*y1�ӫ���?���^�?�%�I�o����a�ō"1[�t
%~�=�˓��(�o3�Xݛ�7Ц�?��wZ�*��W�����|}!&�tPk���C��'tZ�%�慄+/��3B�XXI���5�GȎah(n�"?QK� z���S��:��z}b r��������� �����>���qL���=���3�!*h���l�4 g�̹��	��A���f�5�Qb|������1�dp�^PܴE��pk���>�GL?@���N``�ؙ��&g[^(-`�G��mOp2~oF�A���Х�֝��l�:v���*_ddq�ҟ�dG�`��&��C0��ZқD��+@E�m���P�('A\$\W�y���_�',�$mo��Bj=�u��+2L��oGqq���at�KYa�EH��Q�hѱ�:#Y!��,t��!Nd!���5��!���N|�|�$��Z���q
j� �)Z����S���a�E��P&tgN�����nb��M6s�>G��+�&[6�E`/�}�>����1X�������y�8ɗ�K���W����椵.��@?n=�T7Բ%��O�Ѷ�!�&Y� �=1#7�Y�����D:%���	|����W"�����#ٖdNْ}����M�5n���#nӥ�3���w���͋1�%�Q"C�s͕�,��x�u����E���2F����5�v�O;�]E`I��@��}?XlxV64EB    38f0     c80�0�1A��6�'5�$_�7��}�/�W'��ƃ�/NhҜ%������/&㜳߁�t��ORk��q�+��e�ë�����1�zϊ"!�߅��Dǹ���H^���d@���^F�?=�K|O#E�]׈0�|��A�<����H��p���I�J�=�9wۍmo"h%"���J���Q8Ʈ��A�ffo��Fw��A*�,���6�+VO���^4ƿH!$$O� ��.:�i�,�.iKJb��:$�ti�\�œ�����;�ف%���e������������ݎ���� #���V�##,���'h�6g�a#N �7W}����1=���@Y�)��������4�)M�0�Sff��AV�kF�� GG~aed�y���I{�qdh�T����?���e'ly�����#��0�{��_���J�4�T�� �[ku��n^?h?��`E��Q������Kߝ{}!�KC����k�T}d����G���!�����3^X�U�]��_����{
J	1�^��`Ij�K�5�*��5Nu�b	sf�a-�m,��Q��L�;�vyݺ�#��Rv�?xI���˽�	���	1р�DI]ev4�z��2A����-�B�M���	x?ڶ�A�++M������8��I�����$��䧳�#�w�|�M��J����� �\��Nٹ��vW�\�tߵgu��@���X,ގ+�b8n�w)�L�伛���ؠ�P@���&W΃^��[�m���(!k�k.��]"|Cs�q����N�a���y	#/ �8V���w`�����l��ڒ�beI.�;�N#��ixQ=\h��v��˷��+�t�1��u�h#],�$�]��_���N�Dx%�^:�c8��EE.}���ͯ ��F��" b��s��I�\�L;9l�x~o�^��2I
*�55vz��H3�[�	_x���~�H��0�;�;��uD��y��bJ�c������9꼥^�7a@�;w<]��`E(Ayّ��]\eBD��l�O}�j�g_ i�}ݨ	�t���3���l���B~wPٖE��1��XJ��X�B�ܞO�o�F�~��`����C{�0©�vM;��C���#FU�>U&&C����[�/K	Iʐ��3�[R�;91����!�{~QX�u������
<��=�2)�xd36���PtkOM 
>O����X��<Z����fp)�B�jH奢U��Vriv���wF�ds���v�]I���GL��=a�&�_vf(+���nS��{���~�ıЪ9��~N��ҹ����-}K�C�j�g�׏��Qm� �B���P���N�Z/����&���YU 9��U� C���S!��9����@aS�pu+\�b�5�q�D�Z`4\j!�R!b��.V���?a��'-�%�'*����k��R)�B��y��x1ɻid�ԟ�0k^Ӥ�d8��g��صR*0:�;2���uǷ��ԗ��z��F��G��O�ݑe�Fl����"�9`��{�^�Xn	�v}�>��o�p����
m}����ib#)İ�ACF4����@|C�z��Z�!y� �T����TW魮*/b��[���k� ��t���: u7�z� c]�٠�b�%Sn2 vU��#��S.�2�p
ֿ-aq�!8�t�ϵ�0}��#l�n\�LC�dD���e�3���N�� �����re_����bL"��Y%�	zU���x�����?�ᡫf���F�D�Em�^�Swqj9c�\�T>�?�~�E���c��E��y]���wIu��M'������!*�Gj����@��Y=�V�k�p״�v�D��ɰ�a�� fyXm�'�j�sI���]F@�5ÞRX�Pj�-X���ⅻ�[�I��3����_��EGv�s��v�PC�����ף?P���ۆ5��fy��>�Cz���������-Q�
�t�\�s�|��^Pj:ެ9ZI�
��s�16X�e�p�¶���̓�E���ި����8_aMʾ�1)�6�4��U��U9��~އ�툹�2q�(���i���ݏj����R��x�f�+�__��L�M�ǣ��G�g����4��K*�n�p��@���5�;P��Aꃞ�n�����;][�Hly���2�e
�K�]RRz~mW�.1pD�X�*���w�P��ӿ7�S_q�_��\��N�^>*�q����<��~�jnWs&�3�X`y��A��;V�{�hm�6���SGt���̄n�M�4���_�)��`E*��M�>���<C�琨f<���ԡ�}Je�d�D$��IimF�E� R�l�j��W5[����؍�n1��������~�/[�ԅV./�2�+q�������τ���YoP���3�VsXT��6� �2{O�/��r���$�<,�^��V�_��B��VKޚ�I����o�>w27�@y���x+�
&�����'�"�L�1��630f<��}�$h{�<�mp���UQ�5�����q�fgS�/N�Lvm|k'�}�q�)f?4�a��O�r8�&I�?��G|퀤��E��Ǚ������&��x�H-�@L1A4?��uV�E��6���ΈJ	eK�Ue�k������!�.iY"�G�'��#ݲ�ӻ�o2]����5&'�t�F��q@��{Kfz�pj�:;o�ss����>Ӱ��>H�d�x+M6�z�bu^���3x��Vq\g���4��]�9_I/I���]j����x��
��c�e��;������B_l\1$}N�}���p�2|�A<q���9zc49�x`�)�J"9�X��[B��1?|�&xQ�����2B�<�o�f��7���Z��B{H�S�����%x2R��]A�!A�D��|\�{��ܜ��{r��7r�����Qƀ �w�陽ڮ��?����f�W\�Nunr��k&gTc8�"�V��������|_�-Z�o����5���\��I���4����%��ϲ�W��Q�\vuu�瞇q�7�2Ȏ?x�+&?߷Q�>��\��?59��i!K��G6�v���Wf��I>,o[&���Y��g�x����td"���[k،�-+A�-�C���������Ɍ��
φ��LWwE@�q�90X���.R�%qEf��