XlxV64EB    53dd    1130��|�%��00���9F�,�gQų��2��h11�r�q�摒ھ�vQ���Y��\�Ś�\�9kJG��wb��p�sΔ��|e�u�O�����e��0�U�#y5?���.��] �����C9��Z�z��f�+�
X.9B���U/ll6L����I�����-�`TVnmfԙ	m���͕%zy��gc�C~��Sl�*����m�+�7c.��@<]ʆ�3$�-|�t4�g��.ԱP]��b��� ܹ�F���!�[*�3*�c�W�C^Z�كv�=g�$��Q �?��}���D�侬h�sqN'�8��y�+
2����׏�X�c�������V�4� �C/��T�2�\�{l.Ὠ�ˍ��X|XVkv �a��y��Ϥp�	�¼w�x'��kB��8�2sM�Y�AΗ5�.��)��o�1xM���4v�0���v�����cvʁ����~G
��bZ8�M�լ�&��W:~�b�`Y6����L H����exl3��
������5��?��Ǆb�6�����gd#XA+$vt���U�4�!)?�~��}�k?+k 拏q�HD�E�ۣ�me0����Uv�_��4�a�6��f jHI�ȼ�8C=dj��,�4�;ϹW������u=��wj�rY�f�Z��rٸU��ӄM}��}�=��vUB���~u~o����pfVg��B��!,���v��z�7<��&歡��Roc���Ua9	���
���S悅�>y	�S ޻g�h��bgh��ŉ��^7��Q���lGR�W"�h�����;�l��ɯ��߿���NXiM�����3��ԡ	�����\�i&��-���<%ο-E�����]r�C]�,��g�_��J�z��FUi�*Rd��+	�-K��I(k_�>��	}��PV�PktH1�O0����)y���~��\]a] ���UԳ��SG{��ɘ�R$s�P��X���xe��ߝ!ֱ�-x0_���߮�n�����0,�G���B���r ���&=��v��q.�ǜ���ۜO�����LЄ�TǬ��'��K�@�|�nS� �+>(�����(���W�� ?a�,�𺡱m�����2W�\	���X��)��,"�T��
��M�,* ���F)EYI＞��I���3g�K�Z�����k+C��Qϩg���+�{OdC�H�3�Ҳ�"���
l�e�m5�0�@4��/w궩g�r9��>AH0s���&D�x��r!4T��|�֢�����-��/%A3I�:��-�j�Xg�e��1A�䝍'�P��a�_�c)^]�Sf�����k�f�I���v;�y��ٞM�ͫ9asw}G���"NH޸,����}'s#:��vhZ���B��̄	j�ЄqM�rȣ�^���E(0��y�%�KQλ����vb-�/-97�G���L�
��TvmK�IVr�W����1.Q��X�-��RY�J�U�;�	�s�C��b	�
��T�F�(p�⡚V�I�v�?����.���Kp�؈�,�6�ղ]x�4/�:0@YLh���W8v1aN��G��T��o�C�v�29?�		������(�A�P��9������Z"GW���a�ՎR� n#��(�)����Ǘ��e]D+� ��J0�1�P�_oH�0F|��;� �r�����o�J��L��4T��	�B���jĽ�Se%j��w��T�fG��e�t4x��@�6R�J#R-��%ڦ^���!]�أS�O�������Ih%�����}*�Lu��\竍�8W>fO�
έ�[!���E�~��3\�=�q����������I�����i~�̟���`��Q�p-��iM����h�&�Z���A}��4�K����`pv����4����}mR�[��]>[T1�.�q����C9B,eV;�z��b�N�w�hp�S�4��1��֢��k���h���q��;�(Z�n�ʘ���'v�$���>Eאw���҅����|H�9s�֏�ڠ��?���>0xPE�o�-������Ѝ[�L�{uz�ou��N��f�2�:���$����{ko���e���Cq4?���[WI`�	N������ O8��'�c����2�y�T6eW�V�ey9=����]Bx���˧�>�<�8LN]=z �4�2��'�����D��1fo<*+���1gj���ggY�os⧊�S��$W�P4�Ä,�r^�B�ZJA- �<��8����kc?��­���4,�$b.������������2�Im���qٗ��,�O�� N��&�\;⽓(��F���5�*ڔ�~q1��� ��)t��n���Gy)
��>�������C��TM�E�ح�ޝ�E�+�.��7:W��O�\76Ω�;��z��ϗ��Ei�,w����VœLvF����?דB�0�w�F<y`&JI�y[t:��l��-���!�������ءp�r�3��
�bG�Qr��CRK�r���﫹i��h�az��i�G���#dh��f�T����Ǌ=GT�ȿ�G탵W�+���:���� h�+�ׁ]?ݳʾOk|�v_�������n��p�g�=�+�Qc�>Q���-y�����Q��Tdw,�����6�]��BՍK�
Z�w1 ��y�[l&x��iB�D�FkF���ڻ������&�(�#Ҿ?��[	�<�	*�-��r�Q|L�"<�o� ��6�q�����u�N�dS}��C�Ԇ1�\��,]���MȢx��<z�ԕ���[{ M�ۥ
U�#J�;���Gh�<�["�@��ѡ�i��+|1���C�-�4��5���O�ð.�B:��t��p8 ��^B��_��d�d���հ�e�T�D�Yb�1z��1�Z��%.����&��mt��)��73�D."�0g�Ӏ����m~�}f�=��&�Fت�j�]���J3�vf��J���WO�^��0%��D5�����w����vhS�t2=���ls�@�+G����3��]f:���}+�<���4n����]��[���E.���9��]�C=�r�ڛ�كP�X��F��V�rV2�Dţ�a,��乿�yue^�M;��lo��|%8Gt�Vi�uO�EJ)���3H>!L˾��gx���+�Uji�&	5iLA�خ�s�c��]>C��FO�;�2h��������[�mQ_��x(G�ugn�QZO%��}�3��c�/�9?owDqrٱ�.b]���١�-�����$��Ybߴ��w�`��O-M�W$ԑ`#���T�z��Ļ�0A���>q�4O��v�m��HQ�@���O�:f�*�܈&-�Ŕ8rt䫑"@���'��.�N'�jk�]+�(zQ��;��>�
�V�ٿ��ԣezs|;8@�f�Pշ��:�T���D�e�vt�^��$��u����(
�(C)f_�m��ϛ�;��?�S��/�(���M3���Wٮ�6|�F�~m���(��H�
Q*�����w/`_y/bӸ��V~�Dʕ���IR	���'Ү���*�{%�� V1\T�����$"��V���/|S/�x
_'뇫k�6P����Y�`�u�_�a6KM=��E�|�����eρ�j�-���*�������{2v�Ǳ�����:fb����$����z�[0���5_4m�5E�ċP�7N}�ٟ��uʽ&A+���F7��hVʯ��%ƤF���L=�Xq��K����T+B��Ԁ�N�ח�Âڢ9׆ ������u��v����}�A��[��BL�3���!��,�Q?ړCx��E�էoMy����8f����g8�j�ᔝ���#s!i�;(�>��CN��C�藖�eQ��hc	�Y���40ҙ�"�K��\j<+Qz��||��@��T�	�߉#RQ�A���5��'^�;�1�7'��26d������)xz��w�9����p6��+w����T:���,�guѡ�����E� �-�u��{���&c9��e^�`�_�k���<d�:�S��w��4��)�
%��Já��VF�}6���G���X?j)�z��Mr��o9w���yf���\F9�\��x�<W�ki�`�ףCm��Ip�&0��og�JW���������Bݮ�� �RΏj�l��sV��a(եI�\`0$���V����~�_2[����|$����TP��:k�2�����ݦ% ��r�4+P�,���.�lWe��vVb��o;��X�0�qH�Ž��̊8H��X|>P�T���� ����ŵ>h��brޞ��.�0i8Ǳ�=L�e���G