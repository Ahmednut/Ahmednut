XlxV64EB    5290    1510[�vD%�o�!X��X��n�����+ӟ'���њ�֞���y`*����lc�?c/>`orq]���Ml�$�8�N�`t��H�v��H��!�^��*�w��'�2�Q=+���aL� �Z\܍
*pV�H�,���"'q4����i���Z�����=~�&#GN�Cp�=��:0B�����ES�*% .ֳ�ۈ�+�e-u�}��>{��A���[��Ҋ��Q�=�T��u�4O��B��9;����*J_�CyH�����f�ʑ&�mW@ԗjb�h��֚g	�{�)�̫�\%�s�װQ�a��G=|�Y4k�+�Z�]�v���:�_)��`uR"W���+Մf`�G|ED�����O�u�r�J�kT(#�X0���.��.
�e	�{ƹ�����\��AjmU��%vK~�Nb�
�-���/mF�T�F������K��b�.C��,9�Ғ�H�>�?Xp׭�t�4x"-	Jf7���_~��u��#W�a\I�`3�aHu��*j'�#�hkn�lñ��S��Į�S�T�[W;S�Q4��Ԍ����B�Ιmb^���m�p|��,�S�'��c�4��1��3|j��w'��E?CɞZ=yhQ,ߝ����_R�2ď��.J��o![ #�陊��6��R����iE��RK��2�Ć�Rgu-p�ɥ�����d�G<v�V�;��d�$]i��oh��R.�g/q-�}e6b�`���0�ಁk�?t �;'�xo����]
��Wz!%���k��[!Tj�ha�V�n�݅^;\��=���b��y	� ����>1P��M>H�Q�2;P��! �լ(�E�����p�	kl0� �`�ENPV��秃R�6�K`x�h�:(T�:�JH��>A�!�-��z��ߜ乗
�KƂ�Vlcs�6�+�6����J�Y�*h�_�bXa��}�qd����d�INxس���4�A^��c\]t���ʼ$ ��2R �K'���?{���RB�iF��a����8��m'e!�Rmx��V@3�L��%��^�� &=���gN�ΰ0�֬�%9��� ���F�zB*����T�W ���=��U,�	�G����H �/������Ʒ�=�&�*Fj�j��7�2x͊a"�Y0��*��(��Č��9�]{�T�H 6R���_e����P;�4���Z�G���G!�	Mu�����Յ�l�`�2�0T������Up�L�H��Ac�̫����U���?<?�0H�l	5��N�(��;��w]���&��#Z���l:��H���ݵekc0�u8�s�D�LzI��e���Rb9�.
�z��T]VU�v����dkw����/m�����M��*i��I�R�t�����F��)�|z,��x��]�蘳Qn�	_��|m
 t h�/���Wϼ�V�W�J�9F�t�d�x	1=6�w��1l7�rd�|�cF�ǠR�'#��ú@������W�!)�����5Z���ٲI�0��@~;"X&��r��`��|�4<FQZ��m4�@&M���)����k@�8�@�4	�TOh� B��K���տg	/szY>BqR����J�}�`��D�R�,Q������x2|� ��"%����3�J){"vM���P�UN��z[J��
�v�q����h�6� %vi���J���Q��ť��o�Ѵ$w�f�F���]�a�Z6X�(��vg�tԗ�}�贶��ij�X-������Zξ�GGM׈����4���2��m7Nu�+JMϜ��N��te%��&W���Z>	Mi�%�<5�V����bN
J�A�)��t�����Ű��13�{ij�N��p�]V�6��1���+ GVmF��3&Ly�
�$JHnS�����tU��.;eq�� �n���&��@c�@a�C�ˠs�qī�S�hX��z�lk��]09�v��~��g�zq�t�4ww���i/S׏�P�a-Jю���8�,�I��%�Y��V��wX`t4;X?�zęi?�����or�S
�#;"�떛�_��t$ȴk��Q��z��������&f�<$�~/������=��y7���%���'J���X��y�8#�<Bm�]�g5���7��ӥ!�0�怹W3M�&b���oQta�� 	�
i�@�C���8z|��W��o������iQ�kv����t�y�wk����r����y�u(�S����F��{�%���{c�Vy��D���|�",xi��D��0��[���L�O'�m��Z��bj�Qa�R��F�J�k8��+�^��w��=}����9{U�F�Cxqh9(��y��])��R��Ȕ�/l�b����wFu:��\��o`ȃ�""�e2�M�A�s}�Q����)�Wa3�	�ȯ����*:��d���1ު�{��B�Eh\s3��c�����qՊ.�GS��� 0?��z�vF�a�G��������#��Ρ[A��&�=a��v�΀{�1 �M�%�p��j���W��w��^E$�����7�S4�����io pu/��fg4��ѷB ���=g�i��D(��Js�e�l���NSбe{�O8_��*�% ��]����y� �1 w���t�ɔ��S�-	:J��_�Y��4�2�f�U��K��Y���6[�1���a3���r���s�7Y�l�Le(����G5ĺa��޾�Av�{^����ӑщsN����;,�:�Z_ ���%#Nv�"L_�ל�|s�0��E��� -�4j���.�( ��"�&������{M���B��`�O�#�!�S�~�\��x7\���,�� U��'.D�1Ζv�jڍ�NDFv2Cٌn�yi/��o��x�
!�ٸ�:��K��smɰ�?����NO]��a-sx�26�$�?.���r�k'ʩ�6ζP!`�D���i
� h��$x;XN:-9֡ց���c������֋���?���ܗ	��w�6Zm[�iXyK�����+�� ;z�I58!��ɧG�hjūb=��beD<l>(��IB!b��ȍ��v4��Yq	��^���v��{E##�S�[6�o���݋D�t����S�5��߅�A��a����7��i�ʿ&�SVf��з�Hq؍�K%?N��"5�VN�KW�U���D-��_����+՝�6�Rĸ-1l�9|"��c�E�"��Z�\��zS�~� �PB�BE�V�����잆��e��%��
���ӿ��T6�}$���_i���]�g�C^�n���L%���>UG�T���x\��W��J+aؔE���B����ύx�����T���Ju�jf�c����VZ��]�����0
�k<|a>�})	�W�;,<x��*^���> 	Xa��}�9(s4��Uޘ��I�7!���D`�$����<�JD��|W�������#/e�}G ��l��[�%Y�<S��48���c8�K$�H݉��jB����,Ve�Q3�u���.�+�׉����&���a���[��C����k�`��yXz��!��!���[�|J?O��"���VIU�V�}pC�ܿ�"1���$�OBPC"�fo�	��wA*E	�e�)�Ә3��=M�zd�YN��3�����&mw�L�uCV���ҳ ��`	�������,��A�`3�*�����	�o2g���㓝]{���\_$���=�J%����3��d?OD����'��w�w��A��@pt1�k�=IR�^� `�g�by�o>�H7����Ֆ����Lz��蓽��AB+�	_�ϴ�@N��p(em�9��~fYo��@HҊ���֐�}~�p�ݧO��H�*��=x��;��1Vn����;��g�(��3�K4�9꫃���KBѴ̧KK\'7Z���A�	1N%�LJYC�_(3t:3���T�)�����)��^��rg㛦`��r|W��k2Y��į&�q�^c.��6����`���VO����I�!��XÒ�-\ԌJ^�'ЂϚJ�WN����1*·��g�y��[��-���Y���}]��~K�.��[�m�a�_
�����G��VU�=NI��G9�����im��,�u��nY�r���ߗu�pNYTdkm��(����F0����ݦ������J�&g[��M����Ɇͭ?{������ֻ.Z�S�'L"Z�IEg�h�l~q��Qc(�b>Z�P� V�a�b�
Y�(w�<�~:Ҧ������n����ܔ�O��U5��n�v�ęO4\��g�p���ݍ��͹�ok��i��	 ߘ_c*�H�E� �?�P"�N�의����/E���z��[^���$g��`�e��ULc3�1���0�o��9F�cm˕&�O��� 9�Ni�� neXtԬ7k'r�\�i�����"�3Fp�#���(�T���[Wy�Aq��5�m�WN4�ؾ��ф�`b�8c��+v9q'�w�j�ї	ez1p����!���@>\\r�TpD>O���^���!B��,������+�Z�j��,���f SuT*�����$����i�
{D�\�E#ǾHd��E��,0��c��=ٱ �?�=�.�O�$�T4F��m�v
���}]�T�-��%o�^���eVQ�4���>}g,k�s�G�ޏ]�"�q���P���vE���H7�nV����|���o��eg����1~��U�E�q��ȡ���������d������I����3C
)���a���'�'wd(T��(��*'�Y����8��=�,�&[w3�li|�'}��V=Rr_I������TT��Z�tAC~��cQ�(pM��)ԯ�N
�t��}�W�8��M��ͼLly�)b���$6��eO��o�6n����o�V�i�<��6���ymX$7�5�R��Z�n�ǝC.����RU��F�{H�w����#�m���I�I�������vWs���^��>1�0p0�Vݦ��y��&OQ�-C�>m�ϕaq���m7a���a.��-_����Sys��U���&I�A� ��*z�A� �f�:9�8f��a�O^nY�ۃ0��j*�lh�g�$�l�i/d��n�{=�����
�cN�F�߄�R}3�8kw����#*�+(�ۨ���?x���xs;@Γ�F�U��Uk�C��ܰ7lxf�^F��J���g^&�
ڽ>��3�0Y�9c�a��e:�ùű��p�f�(����E`g�Sѓ
R4