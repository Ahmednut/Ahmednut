XlxV64EB    1b8e     9e0����T�B)��=��V�*���3?.�	�s��
�?�@R�Y�F���&QK���	@��`�䚎�`���o(�.�%=�\�d�H��g�Vג��?�E�&�C#��v��̨�;e�uwGj �l�7׃g�ȠI��	�/5���BX�X�׃26��
w��9�⡂���l"4��ջ��������%����0�Ҧx���֨�c>�����w�����T�*��'� �s�DDq3B��W�u[B��[a!y=&�M�7���S�4��_*��R�����v�����nw�$���Ɗ#νx>��r�+y��	�6��x�)����<Md�]����NT9v/���3R�hͧ�ދg�I�̟X٘��{u	@}Sq%�ͺ������wc.�nr}v�Md;�9b{ͧ�!����5�Yaޒ.�O���E�i�H�JՉ��]�r�;����yB�&N��;7���Ye��'FcOk��J��Y{��.G���1>��ђa�12�	n�z�sW�mNA@�-��TeZ�o�(�"���w�I�Z.2� J�Ǥ	���[�x�zvs�F�&u<�Ս_^Q��q/��I�]�BP��X��aJ�S�l6XAD-߳H�N�������^<�/�7�4-�^T}&n-W���nr[�^���c1|� ^��&��ݺ.V��#��? V,�D:� m�ك��Sh[��|[��%�;�=�u�d���מ-�r�*R
0��;H����"U�o#NF����x櫋5&�!�f��gty���B�8� H�ϼ|˕	6���ÂXh��2ٸ�"��KP�@���ɑg��j0��n�.�LY���P���c<ۓ���
T��\陨���JuB{�������ϻ��}��ޫ�� �h���G{�ܭD�ZŸ��3�����,#������Y6��\����/���0K��5���~8ٯ��g�ǥO,�#Hf5t��)ӡ)�?U�c�qBF�(dȻ'ަa�M �O��Z��	.��}���J��'�sO���~Y��z���>��96	:��{��^@D��B`^�9�E�r���z�,�|��{]��҉,��*~[�U�P
�O3���#T��/9L����	w��$�W���'L?pw����7�A��5S� �V������ p_��Jt�r�r�,M�cq��gR��i�������_��Q��'���0��D!�%n�/���r�[���Dtƨ?�������B�1ϭ�nu�A�:{�[p�_��k4�U�w���2w�҅~��y�U��Ͱ"����tLQ�C�Y_
�?� h4��+$�A��/�#�.�t����&�N9p� �i$��|�Yѽn����H9f	4�q�S�?��a�I#>?��1o��_^��~����N{�h��}���;ۏ�&O�"�s��p6@!���np�(+>
��ќXh���m���.�I���4d�o(9��N�nέK���b��I^g���J$�Y;�W�������	�Z����X�<����'���e��th�F��H���8�-�=�<?��95���D�( D����� �	��A˲1�D>y\��ч~Q������L_�����u)\�H(=���F� j�����A=��<�����K�����;�3���+��������g66�m��@]��&A9`�rIt �\��<���7�g���S���>�q$kֲ���m�McM�b��M��D3d !�"HM�	�,l@��r����1����|C	yeB�»�&�n�I�;�����R�+.��>�0X�:~�E3ke�o�f�R��^��jxE��Qi��k�C�g�o�ǉ
r��'c��1oP
�V <|`���_?�8j� �����
�]ܸl�14�� �(yHq�[�Ƕ�	2�u-���g�)^j�q��h�������5�Q�2�(�+Z.�*��f���az���$����h�p��"j��+��R
sRޱɜ:5��/��䦜;�=��fqL��E�xf�-i�L���Z�E�-���a�:;?$�4�(V6�1��
E)�υ%
���0I�e���oZ����2�{���ǌ���+�BI�{f!�a�_/�0�t��a{�9�
�w��#=OB�$�.�D�
�A�B�wt��@1f�V,����v�4 ^�nrJ����ktG���%�{��}�0����)o����M��O�� FPB觋Tz�߸����|E�b�_v �}:����x�����+.dQ������Ƴ��%�$_�:���h��|BFz7ʽ�������Q��E�b�z=N�_W��-��Ⱦ]$I��2(4b��f���p����|�ƫft�)� ��]m�& 3v+�����L�uo3&����<,g!��c�����nw}�'�H�9z����#��.���>� ���J'�/�rt���D�9�Sml�T���g����m*x���2�V1�rfͼ��(���s��jdQ�&� 