XlxV64EB    517b    1220Y��̥�Fc9!��·���@= ��L)�"������LNQNſ<��KL����P���C"CճYIX�� ��"�p�s�,VA6��j%l/z����2�Đ#Zsr�5��"$��"?�i��a��A���xt�E�;ί�й������2���hx�f_��|�e��P�GuG_¸$R��t���.]��k���gڵ��T0�O<d>�g��k��ݥ�h8��Y�n`�o*'NpJ�K�`r�?p	�M%��N�rϘ!�%�ƀ� �w糼~Ǐ�ke��n[
a�^)��)� ���%3U(ל(�j7i/4)��"H�?���&���)��20��M�V�7�y��8����@�l��e���B1P39K�P�&p��uV����j�Iy&w�8&��8|~Z���-n���/�M�����Ũ�����&�쪠&�4���-S�xp\喥>n�?��i�F�Չ��	���z*�M���* 3e[WU'Z�4f��o���������|�8o����6g/��+����&Χ��Fo���N�?b�p��_cL�*b#��'@���!��u��~l;4eF�u����~k"���E7�c$��*�i(`d8��u,�8��Ǝ���d��0ΘOߟ�k)��ٽv����^����4��v���������k�	0{�������Z��}�=^^@<�l�b�{%]/�L[�§�\�97��q�ep�H�u�IE�[�~)C]�S�ޜ�v�!J�(��bR�P�VI����B�un�M�mug}�O��2��AnZ!�<z��>g���zj~�!�a�������9*j\�r�e��=���y�~��C9��M�b��F�9�m��C,:�W4�]�,��,�L3ӆ �&(�!;�����<��|;t���Hd���V��T����!�A��|�D#V��ТNq�큇㙁Ԑ����7���)���)�U�ȉ]�]O:dgaF.�l�NP�W��� t���bm~�f[�\�ZFB8��99�t2	��a�R���Oܲ3x�p���FF��E�M`�X��6�N�:�-�Q�ǅԜ~� 'u&�6e����A�`�Y$M�� ���\Dn�!h�I>0L��{nǖF��zIĨ>Bo�
}��]$��-d�4B
AL@ըFm�O �B�����P'��+2�BJ��^L�\E�c�,~եl1T�/����x�c������~c�nV�o��=47=���c7������RB�N��PG:� A�0U�ǘn���C1�P{A����Q�A ���2p�5��S�O���#�i���3hl<����N�h�����íB�In<��[�&ԄK�l���K���V�iZMϊX�;��8!0Z"B��,�b����X0xd�I����nq����R�3H�;[��X!�����j�e��#�ˡs�lk�|������,�n�0_"��*A������z�.���rV����+Og���4���ܰ��N��]�!Y�A���ŹL�wJƏwF�b�����V%fn��5��mʷF�	����ٴa�o���k8|��/VX��:������g����5�	���Oqz����s��P����C��F,ݺ�u��F���O���-_B��H� Tc�-G�K��O��6�#^m���J ����b�g~��u�KD���Z��E��˫ʫ�������Z�W�H�fGݾ`�1���^��H�3/�i�QRSc�l��#���@sg�����e���SA��gD�:o2Qu��?"�L'�4?)<v<R$�r~V'��!h��%/�7�	���'�	�Ri���W�-��wE�!m�c5C�'	}Ɗv�%�d+�o]�+�e��C��]�i��`A 嬅	M�"w�!rV�F���i�aM6��'`*��[�d�d����6�g��l%F����cV�m(����X�#�a��a�n�tr��0�p���7!�4P; �,���Y33��a���B-���l;z��n<5���4�z2ֹKu���'��r�I ��O�1�6f��6p$ w�O4/(]{��ͤrq�@+WZ�*�-
������R{ޑS��	�z����en�;�0u�v��)�5=�$a��V�.�jtC "��%��jB&$�������w/q��ٝV�\p��Z9#)�`n�,�$U��E$?�ْ,2[;vV��|��u�"՝��0��A=�#��A���dg�~:sսs\G�
�tE����(���.���\�+�p��t"�=U����s�.��{�"��S�~���+��5�ԫSu�7�C����Akw���+�?�u]U1�X�}x7��2�f�/|R�_�2TP��^@+�����N�Ly�Q�}�e��2�(u��^Agb�&��k��4|�1�Z�@3�.z����b��f2�`F�r�%�g<�Aw��`� x$'�v�����%%��]pG�n#u��������x%0����S4Q��(��U}��FO��X����9�v�oyS��5bE���)wgK &�&��K�Y�"�=<V6��BSVx>�?�ц8�lz����Aܛm�t��[�q`�B��e���������)�:�R������I�����L�V��/ߡ5Q98H<�,v�:�K��u���z
�;%\6r�86}�Ym*�oo�i���)���{�5��uJ���������_{Z��J<��vp	�%{p&&S3ک�����-��~z�1[f������i����"�'�/R]�m�Xnv�8���<�>�M.��hE'?C:4.'�6_)ۗI�c7�L�[;�W�hi�E�����*�����dA҆��gvG��� ���:�a����#�=VP2�N��ې��,+�{.����W��Ơֈ`����7�㓏�j���TEm�w�����O�����&�T~2��@]�za���@@��:��X� Ѱ1S�s;���x;y1�۾(R6P�x����Z�*7A��'�#[����ڣ�/Y�e���Z9�k���a�c��ﺅ�gm��'�A7yM��DAݗ<T ���Z-꽍�/�,��m�^+y��D�3C*D��֋qf���D�B,��oL�_�ǭ-�ׯ�}��6�x�]�����^��b �d鼜�Q���Y\��s��g�V|/p�/)�4!���t�[�&}��2����s�cWNS9�܈��esH�T� �K0eڑ&1���-2W�L��t:���;>��e+�k�v��`X��/	9ęF��R6,��K���������X�\�2a���3m� �J�	:����Tk�4
��	 XR�7���q�UʔKE��94v���]b������ܧO�����d�<�4o�G9΁a�;�+}�AQEo.����8��2��]�^�%�d�;�X\��<�c�ܛ����R�A�c?�	`k�=�AӹT#;5��������Vj��b�0 j�z!����~d,��r�^�D����W�}G���S�t��h��e�|[]>t��ۆ�H�����ы�Jh���C��(���$(#IQ
���?�Ɏ�@�(���ia(��R���vۧ���U��^��ww���E�a<8���lm����^-�ᇓ8�D��e5F�r}�����ެ�XeG4�y�
ޭRe\�t��r"��}��a�{��|�E��萵J���y�TZ=���	\Z��򟪤c�rA���%�3�z�<�*�������՚"t��py[���d5n�c�5�'�v���\��9���	ڄ�	�c�!����(t�WS�X/	o��2�E��w���N�C?	$�[ǝ�ThyռQA��q�Lc��ހ
t gԽ��R�* �qɶ'`���s���{~qz݃c���l_�ND!�Z�C@?.��T���z܀N����jr3�_+3�$[�J�5���0M��(ԁ̇kpdh�3�wۃ���ofj=��j7�~˳ 2&�w�/��|��\�Lk(E��0j��6a<��̿Ո��E'"<���
�W3~k,r T9��9��%��y�%����n�r��݅�ˉ�0��*_�%MXM�s=d3�p0*O�Rx�9���ʪ�ɫ��M�C���L�Ć���������xe�G";A�ac�DO��9����y'�E�HD� /�#x�ή�
��E_!�4E7�h�D�cY"m��~���̏7�8��iDW�_iJ����3A�k(�Z�eNP�z	�ѹ���v��g�5�k�Y��I�'9���R7���M�y���I}���(����	�5�ǞL��Y�6�P@��8ߝvo�f�T�P���?51
ǔ4C�i��̚le��^&��\ߐ�،���7S����&��4WI��ـP� /�Q
[<��o-m0�n�6��Ǝ�J#z�c�9�gGŔ�~V�g�k��C�!@��/\����L��);�?���n�K�=<P��rJ����x�(	)%һ&E�[[��JPB7�Q����f1`�Я�{+R��4���g¼�;A\q���0-�ܼO�[A7PIe��#��s�.��,�<�oP