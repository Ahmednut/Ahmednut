XlxV64EB    4a01    10f0XM���-���n��g*Ɩ9�p�N#a2#a_n/��U'�E!ejrG�'e!>k���rZ?�~��2�ϫ�.F�wSq�%1Xk`��J��(0�J�+�18<Dvql�p��Z��Fp���ߢX4�(8&�B˫�u9�?�-E���1zGE��oJ�@���0�jd�E2�P����5E�S���c�&|������U���.��Y�r6�`��g(5�n8�x�Om��NԘ�6ì�̜��� �80A��C��W���2�X��F#�3*o���)�7���L"���8:�Сiy�c��ݒ�����nj�љhk'�؅����I����t�>�^(��j�y���k�-��	��F��[E"Im�*h�Z�6�Qcf�D��Q���@�|�m,��n��~�:�e
0�*��̍ǌ���io�5��J�oX ��q�,��C�VRd%�"�sqD��Z|��62|�ތ��D�a۞fB��)	�Vk���/��P0P`Pi���H�5���mpD�q�O�ԣھQQ�۝,�cF��ʰ6bH��9��3əy����D��ٕ~$�T�r�O���K
�T�G��/z!���Dp,
+�$
��4����T�$��Vn��)Z�2���e�y��r	M�#l���@�#hn�sd,�P�D��Ҷ��֬���HI�6���l�W��5��� �XȀ;��H�bԳ���¦�X��q1��d̗�.=����_���[�����k�R*i�~^���[dLp&�&�ږ:�O0A�����7�,�{/!_~��p�k�g���q�LuP�K�g����)I�^֋�,���cɲ_%�h!$l�,��t�
 ���t='�A59�;�6�1�Ԇ��1<�,� ox����Ѧ��دqL���QʽS));���#��|�sf�P����R�e&�� x��(�To�e�29�ff���0�����(�����cl�jm֥�@6�JKP��������k�j��l�w����#
���|ix�����{R��[����q��n��~j���/_�W���"Fք���2��!�T qE J{��{�Wi;E��Ts�J���#����d�ۈ��ZZ�H���wt{�\s~�=��u \��z/%h�~���a5<kH�`!=�Y�2߈�_oVH��:��d!�IVH��у��Gw=����!?��{��Ų��%ܖ�s#P�Kz�WM
��Vl�'���ͽ�gX�զ�����~�s�k6���v�qr�a޽5<��Wk��z"�a��x�+8��"#�}��Fr��n�u��}Ct����^�� �#qBY��⨇A:���ͭc'"���4���kQգ񞿵|�ҁ��ŃA)�?R
�{:����9��5*�P")KBL]p R���.���m�[6{oP�X�<sP�ᚳ��@G���uW{���)��#�A�ӲCwU~.�\�����u@9a
�~H=�wJw�%3G��^�)�;|���p�G�����B������+�U�5�ڣ
>�"㢸��#��x�v,5�����2i]$���%|vŸ�j���<���E5vu�Ӹ�b#�ަ6ܨKF����>�� ˃J&�7��ӌd��&�{נ*M��9C����sM��z �E^�y���gk+(�f!�<.v$
*��%Dh?1	���?��� [M��鳎��5|3��mI'�d>_�\��@���Mb��.����}T��6����(����a��_W\�D	WiԐ��-�q~Y@j������Y���4:�T�u�n ���u~��d�Z����O3!��� *�VO��5в�I�z�4�[/4�;��mxe =�Ev��S ��{�m�d2�]/E�d+��=EIߥ�媊��$&�~�G;�DǙ�T�Gml�c��k����b��R����"ؼKB��-��&Ư،͆5�#�.�~M9��ט��`�f�&l?��M��X��uv\M]�'�ԃ�)ƙ��.�g��H�t���7QE��⛏�xh�}�Y�m���,�-�݈G6�l�����T����^WQ.�	���b?SL�R��� 6jV�Y��f�<ob�҅���&2l�#q��4�����D������,�(*�D��� U1�R��,!�M�E˰�E���-�W��r��3�Nn��s�;��ч����ȈP4���`�'B�AfC��Y*O ��[f�X�j ~��>���J�D+�w<�ԡ��&Z�Ћ_((�S�"���ֻ��1i�p���Yjr��b��nAj�$��Vw�hiQ�-`!怔�e`�mO��,<1�nv�9�dV�*�#cc���l@���4�U�������r�~�p�Gn��ԛ�:���k�m��lAk��@ugے�)���S"�����qpT�(u<
�&#�P��{��}���R�'�<�ԮM# ՛���%V!i�A�Øc��N�c�o}�#�r�V5Hm��d�E���U,Ղ��":j%��D�AH�S�/%��-]��!�u�����0?V�!�c
F��s�%�`�Vϗ!����߭���o���N�o>��̺Ѱ#�CN���KN��c�IN�r$��<�����HfEF���Od��k�WO��s$��4p���q&Eqp�v�����ͳ���v�&7yQQEcd[�� ����N=O�%�,i]��aH����Y����>��ҵ�b�[�df�KHQ�"�vI��\#�(��s����A}��h{[\��]��Lܹ!��߰w�$[��`/�w��zHnt�/�E�sp5�������zR&��=���X��
"��#E�3I��yWNlv*�#��ʕ���WMg^G��'�Þ��տ�s'C���!��=H�d�= �mK��7����W�A}���ș��W:+ר�e����M�:�Ja���vt^P������}l���b ����K)$���̳����?I]�۔~b�0����X��Dy���1���H�����3��6U#�^0�W���P{mux��Q�UVդ�~t���a���T2�C�2��ڔ�^*�?�`�MG�+�ǵ�9�t�_��u%,�v}����r��e��n����4A��o�$�	�\�[����t��}����ƛ�`�,�zg7��������o�%)P9"�VZ�iN3�������EL�[�ʈj�
�`�?VX�r�bF��hL����
m�i;���� ���)�W�a�1���Ѻ�>�ٵӕ���ʲ����F����%T��1ـԟT���|Ȧ#�^ f�![��F�]+�(���<�a#M|d�I�$�B��wl�ws�D�'����F�`Mή�M����U��8���*|V��xk�g=�Mj�у=mEpo�� �I��rT3z���4^G9lޤ�oJ>p``�I/B4�ax� �����W��$�p�����[�(���sm��.;*d�)Ԇ��X%j3�u����N�Ԯ�&(�</Q�O\��e�6ފN �U�wdJ���+����J��
�$Na���|����	��<�+����H�Ɯ+8���R��0z˪�)�@�
ף���5�i�J�a)�m�G�GC�`���g�[�B�g���(��?��.D~V^e����%#�z�ҥ�rox�x��p�)BO��э�꓄�k��[Q����;��-���R`~l�n �9�	��>����O+��ַ��t��U�t�$(�%�f�]Y��2�|F�hQpA_	��� м�b�(s�y�YXzvO��=t^�!�m�"���Ou��'V�������G.�$=g3����8��\W�a7�k�vvA,��x-r��V?E���7b��X��t��w�FJCnz:�\��fx�g}���� ��� �)*��X���cz��L��$}�9�KV��LD�rsP�����q���-�V�Q9?}�?�d���F`���X}��|M�X�e����F��$"�P�5(vK����v��(�`�ah]�os*�k9�U�cG�����(:L�W䉎B,b�?ՇvQ��AN4��ӈp��1��卽��B��OA���b��U�CK��6d����#��î�����d1���h�ʯN7�u�D��u#�ʂ�l�����%�	��]��H��%x'����S+H�~�q���Օ[$�~"`��G�l�I:R7Q�D������)��P"��w����jD0c�f�P����<6�+�'����z���>��Z�*� ���!��E�y�8a��V�k�$�ut���j�K{