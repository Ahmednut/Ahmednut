XlxV64EB    15cc     810�|$L\q�!���P���sX���ꂤǍ �=�&+�馯�
G,`�&l�tz*F���k` ��V���2��%	fjM�o�����`��<��v�?���r�~�pKPf�]5㭾O�=��qI���]n�zP�3��9�:9��ڕ�m���[I��N��e�H���h%��b����X	�[��t'��prң(�ZR51`��V��r'=�,^@ĝ����(J#y� B�o_9b��/�/Ѣ�XP�?�ue#8B&
��L�W����>3禀�Q���d����j�� x}u�@fj��bT��CSݯnW�J�6i�Y�����c~����z	M��A�����N�k����:�' C���i�Cm����78�>15�&?�0�P���ʘ�V$��.�C:�d��$3����OG4�i�F� �����G�B�;�-^ZŶ�E�Pο ��a
�/�t"ԟ^�l����L|(��x]�ۮ���Z��Z��d�Z�!ۢo��ј�q5����Aa�2��l>��ӑ��]��Q�P��d:�;��5/�<��	�N�0�h�9Np^��e�in�"0Oƒ�
�.54����.�,Do���e\^��N��!�;}c��>�W���X��_v,�P��i�!�Q���3����y?�5���_t{���q��^����A�ьv=�F�
Ч���0�S�Tu٬n���^BfkT��߉�	XtB��'���S�� r�@�H�1�a:�VÌ���(Bu���¥Dq�:!��ܷL�7�]�3�;Ǐ�������6]�W�m�-��jd�^Ճ��^�y�"5�9��n��ƿZ~?�����:�bUY?9̲���e�}�L�����VGf��(q,5��S#��#��9���~?��	B�P�yH�G(N�\\V�_h���Ui}.�e��S��ö��B�-%q�
$�����×�-Bc^j>Au>�`�>���o��� �-';+%�2�sӰ�m|��ӆri�P���%ɯ N�9��%k-�M3m �݌�W[�>�NQ�~�K�5�]m���ZM�Ƈ�����=��)�~��<4�{�Z|r\Ҵ��9֪y�Am�:��e�Dm0b�8���#�L~���4��U����%�oB�S����2L�#�U�J@32�4��)��|\\h뽚�Ci�o�(����?}P<��g4�>q�m�j�9gN����\�8�q�O��=±�*��w�=�^,	�+�"ど�)�[�V��?���8�6�Yz�][��d)}��ni��Q�𾩵v�	�p1Եe7(tsʆ2/�D0x|�R��9��ĸlǕ_�aB��O���x�씀_�fX4V ���������3F]54�䒠1e�p]~me�Ͽk-�����Or�z]|qM�3���?�Qe�����R�DՊ>R�e@��.��ݠ}�]V�)�T�����T�U@9�l?B�����l�c�O���@�AG��><���gr{�^���b���M�p�f���a�vTp��Z����S��(���,[R���:�������W�������t0KCKon)�e�L^���Dܪz6�VnJo�3,u��5�%�,"b�G���q��?�iT��{���KTj5&Qn ��V��}$fe��x㘠���fx�Umv��դ���{�/+��T�]p8#]M��p؄�;��'a�8�6�M����g�� J�~�{��k�dI�?�
!D|�<��F}�Aȯ�}m����8BќY�h�P��ކp|�i[��_,�{��۳�?ک����{�		���a���S�LԄn�{�o�� �8�j�_hǻ� �;�pЯ�����v�J���X��x.�(iG��.%Mh4��N���S��}�/J1	\L>�s��]ShǷ!b�v0�W���u� �lt1��d�8d�h��	�/w%������o�8#���m8�J����ԉ�w����Ί
l�(�OԟK�����Q���9��q>�>Xi�j�n��<�����z����p��O