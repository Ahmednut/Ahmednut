XlxV64EB    59c9    1410��,�Vi��-�/��ej�[՚@@����Bm���\*�Np�������cv��3��Ĝ颇�E���^���7;��C���;T[�;�z��|���b��
u�[cu�� ��w��𻑽D�{:�)��mv+p!̜���|�Mu�����7�[S啭���������S���|�C��p�`���nޙ�:�L�Gd^���1^d�̑�U���H5�
*�� 8tu*
��V���z�uK�!�Y���{f��5܄���ޗY�%�_о�m�c��h9I����Z{$q���[���`�,�t�{�]n�%5VKj�"sE�j1�����:�H���D>�=�y0��C�5�3���ELrQ�P����Xt$��B'B׉�>O��M����ȫR�ȅ����_I�c_#�kk���Gi&��LM��ʍ�os�gX}\糝�I�@���C��Є�ì�����(�x�����͂����U��G�y�u��;�\AЀz�N�M�#N��`$Z���Q�'�U����c��[y�9�.�ˣ�*���ԣ%o��Ǖ�����X�/M]���.�����G�q8ǒF�U��m�<'��|��<��/�M'+�aa��|���v���<Z"�d�����6���	�d6�Q=���!`�
4�T|����K�\S�V6��핽��z�7A'���:L}SD"�bG��%��O��`��H��{SN�)�>�E��$3df���/�-R�He�=^�ڴ(ƥ�<�G���:B%���u+t�T�v6O���g�Q>1�g	>��$<~��-�����)�����"��(�t��]�c�A��5��e(�}����~a/����烀*@-4�m�L�xd���1�Ң=���e�C�+Mڍ��K�2����:���M�I��0=?y2�G��O(#�j	�X��jM���f^	AT�F>���X/=�����2.�/gO(|���K5�kWi���C����s�޻{$G`��Q��m���o鼄�7No$<R׃H3ũ�?\`�rf��g���� P4�)n��MԈ�)��K� K��z�r���v�S�����὞�F�+�J��Dԗ����������`��|�TU,s?����i�M����.&'B�;��A��,�{G����&�;�%-:�
�q風Hn���|�E#*��>2�~������wPܓ\��������R�-�F1y��5��1>��=�4"�F�4� _ (yf��`?C�^�5Cĝ��t����N������[��i��:>}wp:+��cK�De�!F~���'�?NW�[�ǽ%�� vA~=qG����bn�AIhԳ��N��9��7Q��^?\q�"���xuz�\��\h����kLWin,����R��@��{>>�+�LL
}�DV��HK�a/�e5��'�[�}�8>'V��Ʋ�<2�4G��o��		U\��'8Dd?�x�����zh�6���6��r��֔��`�����T���H^K�z��n$
�v�]o�0�v��������9�({�2GX��.d��G�tmԉ�Ny���/��is ��D��F��A�iI�cz�(:^5�p��zC1��'�)��;A�w�8�-i(6��&���v��f�)��d� �����'�����Eee}6��Y������# 8��×����L�'��{d��Q�CPx�e�=��+�
��f
����vD�Ҩ���WC-no�1%������E��t��M����I��_ �.b׺g-(o�Љ�%|$�j���[vZg�\�6������C�͉��R�������D��WS�!��5�I�c���
�a��4:'|��H�����N�[�&�Wi,�70���9���v�ߵ�ݫ�t0��A����H���<O6����&�p���_����C��>%#N�x�~eQ����l�l�$p�O��K�v�5z=���n;;p���e��V��T���xr���k���x��/��S���=RTw'��M�E�!��&ۦ�m��v�:�A��dm�/�����z�JXR@K�/���.|Y�ɜ|�C�ؓ�\�Ej}�Y$�϶����K����ϣT�gZ�/��6�8&)���q.����u2��*4�&�ɛ&��]W��J�-p�Ox�q��I�F������ �+Hw�����-Df����lE���f�5��>��Glf���|)��l�;��,P��Kϯ��%�f���8|�H��v�|�����8�^JL�iR��"7%p~��MU	\����B��Aqg�!����դtQ�����/\7�pn���w̈́��U�������D�^�DFY.U�F�܍{?��	_{>pk�96`��d�$ ���IoK~Ƕ����*�ͬ���S;~e���G,�XW�a��`C-F���y��G��+&�8.�:���-h� l�K g4��U��q(���g���"���ڿK���iہ9�s���5��3o����u畏$��U����n�9Q��leY�\��A��bK�_�yƚQT���	)��d��ѻ�n7�;I�	7h6���\�1Ʊ�	{��hԑ�)dt)��۝�E���	��z���C�9�a_C���	�$p̻�rԬ4w�hG�W�
����Y��	�'Jf<��4�Bּ�8c�y�H�����؝S�'��-��<
r�/��)8cIC�I��d+Z'ҸEم{�5�HOb����D�Tĩ����W=�ػ� �C���s�҉U�M�u�E6���QQo�
��0l�=tkBZ9�SZ�ْO�RN�7�������O����]�շ�]���0J?�8�տ"�nۄ-Y�c��;�6���J��C)������+� ���歹#�  �8�$�G�&���!NЌ�����m8�չ�� �J0�1ާ�[�6	�E߃�<�#&C����%������G 2b�����+���9���
~�G��	m��1�J�2ˋ?j��=#�0.2L*aj�Lz^q�(Z�Xs�#�L��5�s1Q�\�j�]���￴�H��������bG(��	Glb{^Y>r	�����XM�	�i�?X���z�j
�����S}U�Zإ�r�_� �wxӡ���!yg�s90�Y%|����l�u�3q���}��Kr����<�qvn�Ӵ_\�9Q�	�����ױ�mUUpY��h�����/���L�j� ��"�k5��1����)�g�i����zCx�x�\��S��\V��%}��lͫǭ�)��N�3��u&�#�BE�r�{��ݾ��Q�O��\��5}Kp���d :��WA�t&��[����n����-�L=�S���X��MpU
0���d�o"W�$ýl	�=����h�5�n���i�tT	���싐tn���X�w����b�8Y��a�W6xqۤ��4�F�Ӯ��=[꠪�<� �u�����k<I;�Ƿ�~��1/lv��{�:�����)�(������amԷ����jg �'aδ��Ϗ=,2{V�mu�ᆲ�R�.�d-1��q=�jz�'�`%8�!�E �z!/����e����Gc��zb5ɜYy�|�����ee����^��xChHoI�6�)���=������ ���T®'*�������q�"b���s�W���ʔ>�{�h�_����
���b�UMj���3�O�<J�UT�>� �7���7����ڠ!���Ân�0R'Ͻ��T3�6؇��o��Ɣ�K#Qe,������.�#B)�1�AMZ�򦒌�V���9�7P��֔{�cƜ�� "���ծ}��SLYŭN�Zw~� }�� �L���cUv�m1W�W��wN��y���4Ň�x��%���AM���Ff���3z*U �;4^r�K7�~�tj����[+��
�+�y���&1 �������/�tU/�{=¤�i#cq�I��A��2�J�d?j��o��"�,V��T@8�����8m典�n+4#ۿ���&R�Nz���P/�-�0��ٹ���s�(7kST�ύ�l��ub����ǌ��N7�1�k����G)��s��k�-�B��|ŷ�ZӠTMLΤ�5Ȭ��L���,X6�6L�p��I�9_ʨ0^��E\�X�<(4��1-݄�a�J8H�D^�M9���B�1P��$��.�v���_S|���kWəHS��w����ߩ���у}�{�1���w,����g;�	�K��#D�[㰨y��<&�2��{��`�ɭ���������済�E̝�5y5�����c���급X=���r�i�&���<���KMO����GV��-+�g3���R%�+>��@��/�V�&=��P��C�v��!-�ҠNmq���Ma���+�]���ռZhz�Um�-3Tb��Z��L�(�i��������pʠX��ε�d3�Poiq����g�D��V_f]����r.2,����&'U�пP">[��P��H��12���i�;R�\�RX�V���m@S�W� �#�hfJҲ*�:7o�k��c�[�K��,AἯT`2�)S�Dv��}�^�w|���!�T���q��W�+N��[R�L�`����K� �qB_�R��G�~��(�KkP;%đM��B�'���*��Mb$`�1V��w���<N���$,aZ��Ц{�27(���"�1�n���Bͥ8�Hj^�̞,����<�Mu	Ғ��cǨƱ^��֊�
�|�{�g�0���eyÜ9��$1R<���g�d�Ni���(����Ւ>Y�˼��{�1�a:ȷ�߫B��{���E`�c��Xd�p6}��
��Ba��PbT�b��o{�9�x�ZN��B.�V�?�i^�r	�:~g]YM�ݥHV:&4?�
f�!�r���T�N�3ni��}�+L7�Q��z���fj]��?[���]�Z���;����$�r����/��q�F�-��t�����h�)J���]⾹n `�=	GM=K�M�4����U�r�׶ś0׼q�>U������#(