XlxV64EB    282d     cc0��&�b5m ��Ŧ-�Z���P�䪷��u���S#�#KnP�S\"�`�`hpoO�ѷ���/�swu���h��Vnx���0Z7y�����O3b{�Ƿ[ �Ɯ#�7F9�3"w��\��6~+����k�y)�!~r��g.�,M������]����+W���m1�3�v26׭�T��8"&�|�CC��b;(������j�X�R�f���Q���y�߼X%l9�<mo�ɑQe`��)l?��{	�O�~S�����6?q����� k�鲨^�m�)W�ήOiڷ?�6c����6}�P��h�d��Y�2�޳�ZM�g�g)��v���4�A�i��ʟ��,Y��²f!���ఛ�\�x�<�0h s]<�|إh=��'����uw&Y}.+RuJ7-OQ�
ј��*�<��M�	p ���`#SV�g��s.쫷��p������l���s���-��Z*KH�{!)������$1Y��D��s^��n&/س�V�l9�h���]4;�m	 l��_8(%�q'8��q�&���̈�]�(�rU�<�<��u�>ءd���v�H)Ar���k>=4�ɛ%!�qef��j�i�e�A��{��a�bL�_'p���(a�w8eʂ�O�|���򼺃9�cs�ZB�ⓣvL	�/��l�
�G��ޕk��Z�u�*��T��q�A�x?���/J�4�`�ULq˪���BIN��y�=�!j�%F?��YM9�2 C|��m�g>w�*���*s���MJ�{"��[���U�W�	Y�v�/O���!��dG�����w�p�P�pE���2T��F��at��a%}O#������4�
cb��G�ע@���%@��u�n����8��oA:�b�XRym��	��@2�w|�1k��/��-Z�����z?0�.�����x�P0B�t`�Gn���q]��b�/��<rl��=b�v)�P����"
�Km�i	�����ld�@�L(ǂv���O�	3[Wp̷�әX�3Ɵa�C�3����h��ď��4���G�v㎁��I�v�7�TTVд������4"rC�	iwt�3$�u���������|�	�����8��Ϥ�Y�&� J�D֘���~�E��s���|	��X'�a���!�%��F��H���=#�N�G���~�)Vx	�y����ӓ�㺙������bS2���r:r��|`4�D�/aU��#J̽Q�R��04=�"y�,-��ï�p���
�u���mLX]�`�)݊�� ���M��|X�	�Y,�a� �s����M�]o�&������$yElM�I����)Ap�ᡵ��2������+�Z��`8���9n���խy��{�G����3<�A+�wYo�´�~���w��DA�g�z��75�����0�N_;@���Prz��K�h��̄�v���+�m��a��f)b>�'�,���:P�a�͙ngU\;��}$Q���Y�����Rh�$4�R�ﶱ��3l ��bw돚����n�t��B��/(���u���6�t�T[l����iPS���@��T�\  ��I������H ���[KH�n���M1��;y8�Jj �u Ɗl|�O2�1��ʁǺ1 ,}ZsC[t,D���Z�7`n���d�.�}0�	�
�Rz�Yϝ&`���'Ϥ�2P��0{W�Ɋ4��}L��Y�s���[�+���M��QN�A�%�*sW� s�d���sxt8>�Ò5�����ǳY��`q�i�u�ƹ�O�Du�~��F��g���zz�nL��n����7#��h `iu�8��*��()P��/�W2��Ȳ���b!�iO�ӱ3&
�����э!��u*�m��u�(����2W$4���#�'S��S����ΰP�:t�4�j����kUOH^������Z�7w�5m���C�=�X�M�>�u��q�"�m���[��3��)���6u��@��P���ꆾ�`���k� 9�����r?� �˞�S�\_#??g�L�,e~,�R<w���\g�h���|e@�z"=2HV��Յ���թ�/`?���kK+N�7�"�3�hA�<�,��`,'d�����ڪ+�"6l��#_I*�U�3ƀǩg�F��!�����Y�\�xH�1B���p
W)nQ2��+��>��Զ��*�(��^k0Gv`�K�F�� ��x>z-g�5p��]
���4;pޤسQ^��2i@CS����ԪH��H	���fS>B���S9�����̭ԡ�$V�h7��սi�O�-v�1���Rn����&F��/܂6�������t�l��*��G"+��/��Cq3���j��k�J�����&���<�����k���]�j�e3pڀ��m�լ=�z����N3�j�t>��pi��ْe���������z!���r~�txqLٽd$�wl$�9Fþ̻�r�N1ة]���8x��X��W��3����Cw�@���:����H{�Sb�_���7�]Ĵ@��Z�Ox�-��(b�G�g7uBn��éA�˽W"dDnf� r�a�D7!�Vjy�x���o�YG��>u�T񾭧l�f�cV��KKS�_m���>�Х 2-U{Q7�a�/�v|Sϋ.{�U�p����4M<j��&\|Z�Xj��~� ��i��K�It�q�����r�s���F�t#�$�[��_J�=X"Y����B��F���Mf�a�n��n+�!2d�]\'����՗��
��e�#��k�P�Qq{߈(��Բ�E��p�O",6�`6R���/Sʌ�^�E�����k;̇&A>c�D����<U�b�G񮹦L@ATI��� f p �iۀ�yW40=G.�E<~��5�4@�����|
DI��r}�S8���1ԖJ1spn�8F;Z3h��B��ӌB�Rl�7L�(R|��|�������W�Q�-	�i�as�ZH�AC��:3��@S:3}	��W��.��L��,�z���#�U��Ƕ����6K�Yl����|={w��e�̎z�^o1�QsYi�2K�n ºH���Ϟ��� ��g#0�^�|���������ݠC����Eu�����0pvL~v��_ߔ�.j�vZ�/\��rt�}�s�	�|HK�Z��Vj6E��4g�C*X���ڏ,`1�P��)�F��
��S OP��*�\�4��(�(�>����c)8 ݹ�