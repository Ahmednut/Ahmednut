XlxV64EB    54c2     ff0�ak�@wb)�*A������{*�'������S���s��_~K���bQ�Qz�8Vb� ��,f�����1��p�w�nQl\YF�U�"$a��j*J����ߜHCK�܉��t?���`� �}��CsQ�A��鉄p{PCVg/�8E�[۪�Wv��'���:&���������ht��R�����#�Q���z� V仃��u���:��a\�kj�Y���-f�շ�&`2�<'�5z� 5 ���(��)1��O(:��,��w�f#I*�Y����I�e����)h��[�C������h6�LU�8��2�3ǈz��y0�#���s}�\�ѽ˭�2���2nz�,!e�7�[8��O �_���Ө^7�Z��j�����h=A�x\	�P���<�⢁�9���?[bK$K�?������z�Ut�����l�Fג�7�K�YW�//;�a0�?4�5ٖ��-(�@�޶&�iĩ��$$f��6�q�i�:�s5��.�xY�.����` �o���Ed�q���$�A����]�΅vf,<3��ҕ,z9uM7\�����o�`k���E:(����1'<-��EJ�%gg�vRTZ��?��g,�7�5 �GS�A���2Xã���;�/ �g,�_�Jc�P���H�}~������m��01�¹���!g�V�\���ޫ ����U>�2C2J	(��B���E�U���#����ب��7���R��8��Sm�]�pr ��0����t~[���"��p�=XV�84봘Ì�p��+�bB��N�}�6�s�V��3BO<i	��H��	d�r|�Pn<��sh��z#q�I^@C)1F�Xt��7v�К&��;��{i��%�y����@��ʆk���l<iB���u�U2T�yر���)���z����t�Mw�-V3�'�T��H?��$����'��^X�w�6��4�� �Y>�w?�òF@������dt4�m��۳�G5L�'��ư��1��e�t�i�]���b��%�2��"�!�4��\�R�ozs�MH�ѧ}u1��*�mQ+�נnB��q�'�鵥mz�Yj����EV�:_�O6o�kf����|aE��2ϐ<x��e3�މ���H�3�ݭ���uQ��.��Y5k;_iNX8���͟q�=���@ϟܳ��t��C4|�EU�:�+#X�U�X���!���� K�"�5��-�Pww�me�`	#�)0<%�u.Sʥx��=0,\��ŝ���*V�\Qr��2����Jՙ,�W�L�V�
����!xq�~1��f���\4�������_y ���^�И�?�K"s����ٸ�X��"ҽ� >���3�Pz(��$���꿪�XP���%4�Q�_l�𐠌�'���������R���~B%L�m��'4J2��LA����:�L_��L�6��WpW�D�F�R��{�����^�"}]I�ex^����]'f�|��5q�+��@-]��c�G��@��e�
����t$#�\&b4�bRaFb
��0G	�p�j���ӥ�i嚡W3-��cۻf�5�$�2�1�}q'�3�"x�R���X��d�ń�az���ff�����ON��fu�v�(q�0f&ݭ��A�$P؅�p����:Ob����p7E��5{��N���yQwp`��/��A�PD�Rˀ��}���S�b�b�Q�i�O�f�.�ߘ�V�����S����8o�����+�2����^6� 1�Rj�(�ĥS|bu��9yX��\���q'Lm��%I���e��B.��\��<��lW�`O��PW&�t-"l�\d�[��O\��~#�3"�4X��vy�\���fBn
�O'�� ��g������,���רW�������ۄM����֡��N>3��w�5�`�YB�0<�g��fcF}qGطa��o���a�߬0�V��j?j�U�|V���?k�c�C��CHy��+r���T����t+�mg�����W��h���8NU��_+��p�E�\/(��2�w>�h��3�ǝ-�lj�O���>��IBF�g�,��˹[Q)�Γ����B�-i�@V1J�t)�+G�E�s9t���(��@>��O��!��u.���h֬�w.k�ُO�q�8G����˭�3m>���A"^�+�"y�$��&�a�*�Ge jHѣ`1��V��wy(��n߈�>�K̪���Y�a��?��ۄ����*��|9��O�X�μ��,�#�?X$o��|�s���Pf]�g�����c[����-��h�YZ�m��DW;�����9p��?̃�CT81n+�-�|0�Ss�����H�������� �g<�ANHb���j7#��:�Щc��X��:��~���']�VI�U�ŋ�#�c&�B�i�nK�&3���[�k�f1��
����R0W������"f6��M�oh`!ow) l�Wzcq�)�v��Y���I�~J�uS�<��Ex��
��)l#�Ŵ�C�T��"�΄=�a�/}�W��L/~T�V�3ϘX�R���)�\�]X��UZ�P�g�Pe�r�ׄ)����I�˃Ϟ�V5[�NI��������?%U���b΅ �	���*3MG[�uC��h@��WY̹�r3�*�k|��Fq\�������_�+Q,��-Ug�L�W~��

�1���g���.�ll�:L��|G�=�$�L���8���R�����=�v��������.� ��������b�NDΕ�X���8�8CnH��-�"�h����q\h
u}���)�j��Y���X�/؜��Ǩm3�*C�qС�T�k;e�lO�F��\4��+W�Ӭ������Ͷ���)U�Q$����v��?�n��s��6ߙ����i������,� �(��K:���4-��NZ�i��cm?,���S,�<��Pg��+u~������*F00�Cd��c!�[m�M1IDA#8�M-E����b����P��M9�t�j���y�Q�:xD��>�i���N�oL�;��ܜ�uzD����9�6��uw,C��76��:wΊ����`����?_��a4��u� }���.���g3J���J�C����}?�Ȩ�n+�+!3D�g�%�j���ď�!<�Ɛl� �%{�;C�KmVcv��c�Ԗ$��	�^x��6q	�����]�6�ypz4S�M�����P���)��j��?�����0n�a�6��x$��{o��/���*��[Gb��
GѢo�b�zxq:��$��b8��NP)W|||�)B��b˝P���u��$���-|>M��!o�G�r�FE%R���b@�w���*������s��N�HBZ����E��CC�o�v�F!>5h��iΉV�K���P���x�Ó�H^���u���;^,�	���2�tr>r����`��-�k0܍���N`��������ys�#�'��{E�xO��E�W�F8��Xm�7�`[��n�� 9ec�b���;�	�}�8�'+mpײǓRܤV?�섲���Qxf�v4�$�ǲ�?F
Z��5���7L�@��W��O�xvS��J�ၴ���K����l~�&��t����x��܍�W^\��m���6&C]��uD�A}����h���ۏdQcE� q>=X�M+�ue���w�ER��V�:�� �:x�F��`uE��n���Q�N�l�����J@늁1��r,�5h �$���}�P�U�[���QY�HP���p�FS9>4�rt�m��gM�Q���jLH�u���-0��A{�dO	�+>�&wP�SB������{��VGwT��49��k�p@�5�Zc��G%C��b.IQx�h�S����Z�2kR��Y�#R��ƍ�U�-�̦!�O��7�v�ܿ��Zc]��4�BgN����.?�)>в��GH�@Y�\q��խ/�)��:"3���K���g1%Z�b��r