XlxV64EB    8c64    1530����d���?/M$`���8T��E����dzG�65�mv\w^o`t˕@�~��\�۝h��{��э�v�U��Z�/��)e<0�g�����z)C��E9����p%>7��v�k[�v�b%�/r%���������*DX� 㸗�&�g	��}��b�XO��s����	؅~�+��Ͱ-�g����z,�XQmo���
��3�p����{�*����L��iw�!ͭ(����MP�!�z(lک)X�~��d3�䢚`���f�-��{v6O_��/���Z�>�5z���K�_�+Zf����B岖;�d���旬��dcv&g9��%�Vz5���z)��>KBb�5u1
&k#sm(��w�]+���H��b�PcO;����ـ�;����߳�w0�<����l�"m$`&v�0���G�$�B*q0�-�3�l�k.�/�"U&�C�ު	��(!��K&`�_�)�Dۈ����W
зS���� Q@"�g1��B�@�l��1+��/��
y��.��ȡQ�o�I�cM��e�u����̢/`��'� r��

(�A�ޅ��"sp-蕣������i*
�$*����n��_.a�!h����k�R�a��`+��q����#����mH�Q%��v��i6g�Nn��ԓ��"�=7@WR�������-��:�Ha\�
s(N��a23�d��DR7��i��:=״0Iz���8k>�#�\i�[�g�&cP�}��f��* pY���>�Q*H`]\~�Pp��h�r���L��v��Iq����I����>��Z�P[`�x�l���+۫�#F��z���9n���l��BZ��7���#$"(���R*���[�3�-�_|
�YZ��˚�ꏡ�gR�^�k�<{�3�ܙ���6�pӜ�& ��1�y�p��c"�m��^B�۰u����d[~�
+D���K�Tos�;�����|*�u���3�,#=O?�ֶ;f2��P#s-�ɀ�H [X�{4U�`�h?(��\�/Z��_N~�fjx�c}C�dB��$Nk�P�t�B��	AӱW�\ԕ	��l��vK�2��8%��[p�EGQy�+;��>&�~m���dL�\�L.�7������$�/dI�7���W�:)�W����H�ӟ���Ds�������9"s�c��T@3����`�G4Vn���X8܊8��1Z�X�X��N�*��ؐ�|���&z�� 1pГD���q��遘�*��:}Ma=U��e4o�n���j �
��z�A&�����ӧ��v��1?�����K�yɼ������N�
�#f��� `r����^ #7Gz�,�4�aK���SbjRV��u4?uߪ0�gGU`�}�2�����Oh�0`���"ꀬ��� D%�0��)����r�.��_r��U�6�����X�e%Ó �(��ö|���	�\�4Wd�*���jVu7k�P�z����9���D1��-�`�;�%)�t���xb���	b:�'�{5_��Q����H��������X�F�:-cǆK��05M��[
$)�y��������@����+=���j"<��?"�]�x�~�[&f|�4?��la��k)x���KP�Xs&	(���E�����ϒ�J�vBj)h`2c[�9p����;�ъWA�(&ǈ���Ҟ��ƍ�9��>ɘ�ȸ!��9:�*��kXI�t=��aaoFj�I�|�k�#pi��> �dyP�b}�{⤰�U��6�'6�QċX,S<�[���r��tJ��Yj>\��49'�O�p���u�<��������
�@KJ ��y[�r:��sfl��#����$��\��Гӈ��l��++���>J�X������Jw
�n�{w�ɜ���""�oM�_�Gǻ��@�BG�RD	��/��>���U��S�Ŵ� �x9� yw�U��]���!מ]R������b��k8��v�	k�G�0��{��":m89cHe���KUzU1����
��o�I�o܅yC�ȼ�i�yB��\N�*S�[s#k��K �T�AN�F�f�����2cg��'�mn9�.��rY��SSZ��1��`�h��BO�������n�8���8d�wK�Z��v.~�=*jN"���cl昲�r� j¿�>20t�B�o��L�ǭ�a&怚$f�?4�߯���2k�sR��s6�ڠ4B�����M���DrJ�Hc/e��{��������N�J��P$b?���)���G��]p�V�|;���%?.��R�s�Wn(��>�S�������_;�}Gs��b�/w�?���o^K"��LP����o�67\X��R )Q��r#]+������H��a�WUT�t�0�O�X��\l�WH	1T}�����TJ6�9�:΢�b��k�m�_����E�N6�ޢ,1&g���w��� �/	3��G�<�0m��8���ቭ`�!:)�Ѩ�>��G �g.��*�8�g�P�ا�����)�u3>n����bwL��d@�a׵d��1\�?�d[W���7T�� �>�oά
Y칢DpN�!J*�
�-	�����e	:]���~p��_�"!v߆�'(��dio,<�8=�aQ.A|���*���>�`b8���z����z�V������i]�,VP�m�2{ܲ9���cDE?{��,U������ �b��07v�8��^�^=���7�Ug�&��R� �wxl�֒	{4��]�/	H�$�t�~�1#�E.'󞩞��$v]���Q��!A8�a��㪕�I~�M�W�z���|���k��UB�2P��[� Z`kQ��z�h����p#��ՠ�����z��B����-�nqG~֌�	{&-ՠ]�
̽[?qCD%��9���3S$DE\�7���(�lS���P]�a�t#�`}[��T$t�|����F����̗G�^��{6�zR��A�N���U#�!��� '��Q�Y�HN]:��6�@�W[�MLJ�w��6E�������F�5�2���fc�������&#��=2����m_�ʜK0M7{	D"�!ꬅ#H�^|��0��L[[O��O���9
�H̭�S��\ơkT���Od �}���)�ӨQ2w�(Tm5y�
�շ��Jw��#��wu�/��E� ��__�pb�5s�[�D���� ��P��*Ѳ��_F�5�����@�o��Ki����ir���bk�;C4*�(��畸Y8|:ص�Ɇq�����T������ӵ���[�WA��}#m���Ծ���� ""7�J��ܗ����1�iGk���n%m:Ŵ&��!B�`<����F4	�nGckPy�i��#d�=���~�n�=�T^�Cs�uS����'Y�{��e���79�2^*{.aآ�6��+l��坑k��z�AS����U�+��X���ҖY|Cj���T��ō�$�f6���UCKz��|A�����z��:K��xYQdڶ&+�g���f�z�T��Я7���P�ϢA��E%�h*�������|$��<���w�a��l5HHԕ�f���
co00�u�]���gC.��M��r5D�8׉hcjK�g��'Z�q�����C�'���e�:Ɖ,ё���X��ߩ�$z�&��M)��/�%UT
 ���`���;I���6d'�)�Z'��t��4ΕP�Zˏ��JԄ3�{E(��$�J. /�0u�˸fFDa�C'�՞ѽ([���x�"�i�{��ٮH����~G�m�\)]�F7���L�s�N��(�t�������{X��1���S���*�V��T�'�fW:�dW{�����������(yv��J�t�e[б�F;��As����2��'C �F�x�B�^"Z%�ݔz�p��-5��(�g;q �n>ZD�== ݯt��j8��tT��Aap�H�M7[�x�2zv'��g��o��k1n`� ��F\�2�4
e��N��^� � $�R�����Hjn����=�r��4l]pN�k�+��J���'�����^�����W\CM�C�E����:�!�S{yD8�JFcND-��3�SmKWh�V5�������Ц���X��3ܼ�v��&�Qg��/.��a�%�
D�%I�骄cH�,%r9C'�wj�Au�3X#��GT���I8�s��8��$n���1{k(�\�d/�L$�N���-���{_ą�9�;�B���lt�!@�>�\�EU�Z��W٪����5�W9!a�|`|�D9��;���q�ۤ��fM�������l�͕㨎�,��qߞgi��i��>񢋆���W�o_�#�~Ag$Ǘ�J��Bq.�ً�o���Z�H�[�Zn�lfi��v�+K���̞����ԁN�o�,���kg�(4y�����9dw���1�Z��N�.�z#dhD�%�c2TS`��2w��9v������B��Y����8���5���Y�ZQ�s�c�r�J���n7j�¯�����g-s����c����7�4u�Z�>,�k��.��T�e�m�o�7E\�+�&<e�_-�4�8�Zl�n��P����ĊA���.�Α�̈� ��F�)�J�٬���l���R@���a/�6�)|;��f�L4Ҭ|���(�7tr��_*���!�Y2�'0XT�a�I�X����+���G��vʶ1B̏������ѻPFΜ�v�V>)���c�@�����۾r| �&��}��n7C�ڊ�Ɖ0�2����nM憾��Mk�cp�d�k
�F�6�l��Ё���t]Ѹ���
�����d����Sc��{��J\꛱/��8w���v�����I� �@��v�50~��Q��H�am�#��P�ڗ=[!�e5�Y�V�ʔ��Ƨ�p3��"d��CƳ�u�i%h�%�vP�ƺ42A[+�U�iH�YI�q�-�6�u�L�w�Sv�>ʻT��.0��@�WZ�=�$Ȟ�M(����9�����N╱����:����聥p���F��[N�Ű�2g�3ڪ�]�fT��O��%�1c\��}�dUtW�sex����XЁF?ok��������7��Ic��n&���/������Za�@�����w��a)Õ��z�2�w?���|!_�6��pǶ�~�f*�5�xh/�4�n��Qj�!)?�m	��C�"�&X-����[ܨ9{����
'i	�:�tXhL�P����/�W)m\4j�6��#��9�i%Q��p��xƾyd�y��yV��y���x��c���ez��n���nHW�@%���~*�>=v�. ���+���y�G����hB�*� ��g