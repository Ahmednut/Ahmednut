XlxV64EB    3816     fb0���{���s>�"2B����z�i��`��yj3���눐�o��?W���aV��B�1zm�i��.;c� �F��"'�d��#<>��Vl�����������+`\X@1�l��<�N9C�݄�����=tXo�d���̙�YԂ��ui�Z��`���9t�;w��C�Qd�pyv�f����X}�� v��,������Ђ'J��y�&JB��c2���e�K>�gZ>���֏�uAW:��3D�!4��I�l��%Ҝe<
#h��Ɵ-���.��|����_�`�������86	�~H��u�-�ej I����U0�����c�#�C��GO���X����6หo�"��"���>���%�"y.}h����<m(�e�g%Կ��t��pf�&����QP�z��)���S��#f��
r�ڼ���)�l��_���q�A�zX�mb����~�+��R��kų�C�E�g�C�X�X���>L��fF�̱������=��l-��3b4O�.cu�.�0�a�E>�ń7#���C�˜*{�ޱ�Dd(,��~ċ=����,f�pCh�Zp���a>
v0!�D�ˍ�|��`������Jn�gD3���b�UZ�Y�����7��c�~�e�[l�f�����A�����0�J*���B����|�>��%���N%����6��
T�MF�!��%:2ڃ �vU���!H��:O��s�$��&������#�Rw�2Z.	�2a*�u`z!�M�A��W[��݂]�x�J��#�2���s6-��&���dJ��	%N�ab�H5��S)u��p��f�JЙ�jq��0����M��B���`J�Y�z��.�t����$;
���?��Ś���=uJ�<(���!z�C}�X#v������)<�|�3i�y��C\�t��c5 �d�z�ڕ~������
�S#:'�Qz	����A�ȕ�(�����.�=|\��$��-7V�:Q��i�3���Š$�Z5�˄1�5w�0pHݾ���ԞH��Y�[:C�d*����m�� �1{q��K�2�^E��[\�
��7H��;[��~���+"d)P�Y�>u&u�+1��tHn�y;oխ����P�p�n= ��r4N�|^�cPZ�}[ב^@��\;�e�P�ˬ�k�D�f���Y�e��I��}V�Җ���8��~{@�~�������N7��8	���Pk�r��C���g��=�f�}<4�-�o����\)��2�v�۔�����8����(lK�晇�Q�͎��ua��1T��;r�,�����T<��;Wy��ZF��I8�:�k�`�[HE���'a�V�R�1�r���M�!����޷)P��מ]�������|���8�%�j�	u�;�)�_ڨ�v��0��J�	�.�4�?1k���0V��Wi;���o�G+BfpX�X�ht�P�E�M0/�Է2�Ӡn�8�Q��RCo� �%e\y��Ws�VY7�e�Q�:��;	���|`�G�L�nl�|%^J����m�H�;��:��}E�0e�[�q�ڬE��2)#�3�&�y\�#�!��5���WT�g�@4��<b^A��HV;���'�+����8�7�PI��:O�F����Ki��4s r(���#s�6����^v��������%@N 8����a��$O�����	�7�`B�
��ܥ���&ǘ�m��E�a�x,�&�p ����Q/I� �7�?W� �`�>ΰ�C`~[SsPh�Y��p=+_���� q&/�P5�.��9o]aA�q,_o�W�=-�U_+_]C�D�E>����;��ĭ�4-�̀�^�Q?k��j�*L$b�CR5m?4��;��&�t.�~xr"�j��ZƩ���o�J�徔eS����Br���l��W���!W���l�R#�f�7�����
h[ǿF�R�C%PA�.�VTP(�����s�_���A���[��,hV��Nj
,�Y�_̴YҠ�����v5�/�C0�U=��z�`��3�� =ߑQhbg3��Z;8�(��m�@�5�T��Q(���(K���ԅ����CD��aoa�bK-��䨡�N>7�����U��E�^H-L\�X��6��Q��8~�`dۣg"���m��4a�;�o3��z|��{�⵭ʉ�n�TM'��v+���Kh>�?-!�r�E޼��tPY��e򉋐j޴'�%�_�}8f�Q!Ha�������8�_*�	�@�5d&x�o�ݰ�wV%oWȔ�Ʌ&�k�!~��X��/�D�x�K?�N�%�_,�F�ӂ�W�wr��%�Y0��n>Ȁ��2�'�@>333%��,F� m=<�.Hm D
xażK���Rx=XE/�� �� ��ȓ�rej�0��br�93�1�L���Ódp/����3���_��,�e��0I�W��Z<c�d"h�}O���o��%���i�	*W7"i���GH6S[̀&8�< ��@u���G��o���XX�M�~��/�F��}��u��[���`+�����f�0	w[ŝ����xE�\lzk\hci[��NԞV��M%�[�`/����d�@�;�&DN�|�sf�tɬ*2���i�
D�V��V5��H�J�d$3�w��U��p��G�+bw�ļcH�k�{��Qe��[��
���/��բem�\k�ZD��q����>�e�l��?g��ۑ�V>�s��WE�P{��H���-`V��*s��r)ʍUKYT�N���YnԐ$�0q����U���v�5��\�K��(򚛫��T�zf
��5�Ԩ-�s��*�*I�b��e�f|< jڋA4s]nX�/����!�>���V���1��SG`�q�;>�U�GD<4j/�h�;9�E� �xo��U���o|���.�5�dTȯV�_��~��>Vw{Xs9�4D��@BN�%
�}�e~�<��A=f�!��B� �_�������&�)�G�����	&ꗭ/I_��]`t�ro�������`!����"5��!��.��] me�A�z�#hM��׼PH���}�"	}S��A�GsB�O���������ߦ@VZ��TC�Q=$v��TD�R���f/�+(���F�*c�@�Ra�x��z��"y�o�,ˇwӛ���?75TdRT��/��[��%�v��@=�Q�>BJ�N����Ӈȉ�d�!n���ws5�/Q"(P?�FT��>��PU�"��JK��p�FlN�����\+Z(#@����:x�� �$��TI�y��8H+�U����۪�{/�U@M������g�N����l����	�����[=�*m��~+�����l�
j�A$��_����-m� W���
�j陗Ċx��~m����sxhT�8u��V�nIu��7K�� m����>[���_̜�+�\��u{T��:���w�U%Z�X#x�����Sw�2�?����03��-?��A����蕮<B����j[^#��t>o�给����5���LL�VL$s�0�@#�ʑ��Ǝ2�#̵}�͑p�Z� /{C�)�*5ueY����11D�0$��c���i��Z6�/X���Q���׬wo����R��?�n��'+�ofN������h|��1F�ʹ�c�D���з�C�J44�F��!��s�SxyNɝ���>"`��Y���Qф��^2����u~����pZ��9��h����@K� Yf^���~�x2:q�h&Ξ�P ��(,܊R���@q1��J��ֺ}S3U�����F2"/�ܡ6�-ێs�<rr�^�Vy�=.��Y�~�uOq}DQV��{<;;�~�V���'H�(�ɋB�yڑ�uz��J|���׃�"g���7�� ��|خR�A�)&*Ƀ*�����P{�