XlxV64EB    8a37    1890�~���)�k�<���H�G����<�ލ�Њ^h:�*U��
�4�%#ސ,��3oa����ZW�l���$� ��ή��5P��)� �xB��ց��5I���i���;��X8̶�*��P�kǑ.��Yхc�;��^��4�'�1�mc����e�T��]��3i�����ioV�Ok:_�u�C���@����>5�^̪������:+�dG����fI3�����yBmi@9��PݏZ�β4��B�w7���͙��$�d��:�3~���Z���d	E��US�
��|���-6��{��E���&h��і��qV]������e�A�ֆi�:7�9�����w��	v/�f8蛱�u��m]���N/��o7�$7���&�t�h�K�V�x4F_ 
�g]aU����������ևE-���{�!}]��mGx�U����,�@��	�x�d�_N���4LvU��<A�tT���__1�Gj"	
/�|��z�{�r\���D7�/k��1�_����r�+	�~�n� ���@�[�G���+UL�kz�l�(w�Q�mF��͘�[��1��,8WA�oC;���h��"�I��4�����*�
)�O��'+f�
�3�J�g����ٶ�V���`� ��m�}h�ٵ�G|u��T��OL��~�m;jZt9�����r��ֵ՚��@�\�4�k�{��]�cA���M��?:��R�cJǱp��R��맣-�wX���z����G�޾.w���x��q�Q��8Р�t���A��1����	�z��{��_Kq-ό��K+�5=�qr4�9��ym9©��Ro�ْ���v{?�!�����8,�|���Ud��3�����I��A���C�z��ֶ���:�{��d���%e�"��[��5!Wq��#��~�Ѳ��6��hj+�
Z36H�Ҩ��K��zT����z�\�������~���xӸƨ��^�&l�N�[����_����c��p|�tM�o����V-ˋؑ wH��p)���0���,d@�rez���>�lm���#���y\��H����a�m���������ux�����1��x�t��(��B�%��_�
%5Y~�o���ˈ5���4�?�q+��� ?��QY�s:���M�SLDz��;+赠"D����i�iM��!j�	 �R ��_�	3��]��蔏ϫWݎ�8�\���7�.��M�����;�b���1鱸3��??U��,�e����{���fr�C[���-���4�y�i��G����og��n�x���;�DzM|#$��ƅG�l�4�y��io&�v-�虡��� ����O��ʕm�Rw#�"�]rx_�0�?�.|�kS�Kbw�{r�j�d��0�C�A;W��g��h�݇�/f�%��x"
���/s���������9����9��ly�9NBr%�T�kn��c1��!�줱���^�@�
�Hm����<���y2
=��o�(�����,����C���m0.Ε5�Oĭ��C�=2�k��tlV��^}cLa��]>� ��ɢ��[�_f�8�s^+���%�gVJ_��hq�����9�V�T9�k俅"�j�����Z��Ӭj"UVF�!
90�P�p���u��QJY�����
fF���x1h��2M���<)��|rXf"��� >��m��	Y`#.}��N���.>&[��$��^'��2
�Hz�y?O������~��ˬ��A��)�b�u�8� y�tT��;�0�~X�ve�ԏ<';�s�[��Eo3! �Jh�c�D�bN-� L��]]��<$�����JU�Sh|T��ڮ�M|�c�}G ~,~����YBJ=iM��/�;����7�}�XF�hM�pN߆$Ρ���,�sL�M�
���K�
���Gn�����������I�:
�VC��}q�ᘛwdM����f�" ����"ߝ�&�a�_�n�נ��~b����8��I׾��{��_��$��ˌIoq!��~?N��0p؃�`I���zj�N~4#~�]CvV=���}Sr�����+�H�
��q�b���L$���E�������M6Z����<7�F�(�3V4�pXQ����Fw��&���W��/軩x�=���׀�lh�x���&?t�����j@�0��=e��#E�$�����m�~�U��Q�I	/%����uA����AǱ}
�.?p`\k�PGm���ףJ"l�tM����5��� �nɳ���~@hB�XX�飸-Ը� �9Ek���3+�����O�؜ú�g���\����IL��o�.��v}�F[m��^k\lϭ�^���x�P���_&���_�|2=(�7��nl)���Ѓ(0�h��I�!�@�X����'���[꡾S��cل�"��|4��fq$�[ jƾpy�Rp����*<*�i��a�E�^]���L�������$aZ��٢�0ѩ����l���Cѱ����88Gx}{*	q�����qx&3&᱙q�8/X _d��*�X3~M�I�Scjѹ�o�A���Miz��ǂA3���7ӭ�P�I����jؘ��\�����T~�忴:8_�6�ir*l=��|V H9����1}!H��u0l8z�����/�������A%��
�*�J�)$M+g��\�쑹�rV�܏j(71Rg��B.$��?O�e�p�̅�mC넪�Y�/�	�X�)a�%��̛�ߋ�o.�
U������_�Y�����݄)��i@�&�	����M#Xt\,g��RF�k��%�
R-2�_��"8��r�� C�}]���C��u�J���ko_�.�P6�?:u��EO,�I�Q^)l����4u*�tR^X�ݰۅ�5\�>��%�h
O(��j�w�y.��[���L�Hb|���ĕ6��`���ʭ4�E���Т8/����!��� K�j����:�� =�󚧼����O�2�e�8���9j��'����$���q����{.��t,�@2e���QLt��'�3�(}gl�1Qe�E���˨hx%��m%]1���u��& ��^�\j�Q���Ջ�=I�����rJ�D*�V"NM4��*���:�T��S�u��+s����\��;��!�r�"^V���N�g��Ñ[GUU:8��a�6E\�~2e��9W�h��M��<����K{%�	(�&��,��E�f{�@��ļ&fM�=:
\��Ӏ��yִ�����7ܼG��Y�v�̕.��Yli{� �#;w����վ���{�a*П���w7ǀ~$�a�6,�J��'��`3��ҕ�h�jz�I��K&����5_7�0o/}���kb�`:P��c��	{���M�����֫EC�3��5o/�6�O3f�*;<���g�/�|����2>hw���&����|��n�!���x:UZ�s�|� �Ur�K&�/� �~�Cc�2Ԃ\���d`�wk;���8=�L;J`&j��'�w�8|d�5T��z���!���F���ۦF�(8l�K@f豄�Ȁ8�<���ˋ(Ѿ�\���m�X�i�X�qRv�m�1G>Cǘ{�װ��7��l?��y8�2�]B����L�ѱ���j�|�ޘ�L�'�g��b�8��<�"�e3����ϼZ0�H6�=�f���9�K���\~�lg�G¼��N%�e��1A��g)���N�A>ߴ�t�%uYP6��W3(K�����b�Vº�T�O�fԠ���h%-�-'��Z��a�"���:Rg��1!��1ۅ����.iJ�&�$��LY_8q���V��򇏛�b�uX�m �yl�9($(z�>��r98<���x
a�v,
s� J�:6��J�'ŗ!=J��y �Go�[�LH��E- �z�%���9B�3<�$����%(�nc��m�]�����2]�r�!鐎?`�C]�E���]*�y7S�*�kNUK��:�5�=}_gv8�u�G���m�ٷ�^�X�1�n��~�j��n��gM}�����,9�M�0m�R�[�g���QB �c��f���ž�r�f2�����������E9ݢK��~Jr�����&��Ӓ�a�Z�s5�\g��҅�,A䔢�a��ʄ�Oa��9���w<��B��"��&D�|�BSk�� ���A7�
�i�.�b���s"�^""��^J1g`�ab��sh��
��"�8�{^�t^��f���k(x��_M�{;'�טםP)��L,�9�a�{,e|V�
�m�T�_G8�0oI{�iq�b�%���������,��r��Pgbs��M?8�_�n��Qc.ʌ�7�UL�.<�Q��l��;��4 �A�$E<�u���녣'By�
�L4�<Mf�ą���b���8E���ɒ*��P��b�v	��U��r�:����kh�ƭ��$Rp[ޑ�7���Owձ"���V���B��9�y�6`�F��Vu��P�)M�F�{�&Vr�|���I@ā<���z���t<�M��Z���`W�&\����|�D8����$�%�,\¼��0�AUr�y0l��6g=�O�,�l��W� ���������d��C���qH��2_��S�Q��ʡ��C�ʲ��kI�@���-��J�%�>���.:ӱ��S��?��~UyE��A��%�[��M_v����7|��/r�����0���|83�[2��}l@&(��e1S���(���8�"�OJ1��0���e���]R�pܻ�(О���4f{���xk��1�5�Qv��<�vع�cV��v��5��⯸��eP�Y�����s^S�x�="��ԡ�mT����2��5�����>uҩ;zA=��.�����}�H$3��S�#�����
���!�J�z�m������F�����V�����1'q k�V��P��9_E���uf����6_��_���U����冧��������aRO�$X�d"�O�p����>�k��)4	�rFt��*�$��I�՞&D=m#Q�P[�G^iR*)�a�a2wꆔ�?����ӆ˶L2&<�Fu��8cJut�-i����{dB���g��]�9% beS�L*EƌU�#zX{���^�/��$�3=Sc��{�`���p�ڿS���#�t��ذ�b�AI�z��v,����\ܲG��\�a+ ��U���6�fi-w�U���ߺ�:�yt��KX�5i�^�� |ª����5K���Dp6�mh=�~��À7\���K������bY����<���-�a{:���ш�FI�[���X��d��P��Yh�(wtk�8�l72��m������{��j����W<�I��ex?��F�D���W��~x	��{�,�mfd]�rβRG�ZU��	�P��À����R-�#���Е�D��}��wY\�r�a�v5��F�k2��Q���	l�)�����@J�.Z�ag��5
1٨ nl,,����=9�w_Cl���WV�Y���l�^�Jl���Ԏ�L�����lo���;����3ݦ�v��c\��	������H�!u�e�ˁ;�����j{o�+�uMfq�,\�����.���roVF���������.}Nm0���LPY��������e�䕊� t�dQVW���@�=` ��H#��u���ד98��G�=P0�;*���в
	j��k�q����VK���-Zp��CcE�RR�m�-.�
���A���9���c�&2��ʟ���� QgI '"����.N9��(p��y���l��, 䲎�!	u5�������Q±�ԙ��Y��]^ͨ�V>s� ���EfٴJ:��	�8H�����YB+֡Xz��^H:6�7n�F �GBn��-��Q�L7�0p~7��)�~�J� xe�V�ٛB���{��������Kx�ep J�h�@%$8��ǒ��x�~���YPYn�(:�1��̈U�����.��.�W�����x� u~T�X��9�3�0����x@1��9�'vX?�PZ��H7�E��	�+yI�cF�2&�֔-yE�"�p����	c1g̲RjLr�۫׶���Ks'�>3��\�b%̥��߀f0��(F@�5�3O> �8���_Q<��C