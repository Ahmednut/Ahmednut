XlxV64EB    fa00    2d40՜��'���L�N���i$��P�v��1R�zW����7��p�]��b;�΋��>���v�E���$�Ϝ���e��&ú��>M~�J�#&)iws��4`��4㒈K�چף�Ay�VF�-�I{A�:=RY�
�����Rv`v�o�`�k�a�ܚ 3�(��6�.W �߷��a4jnM��bB�����3O��GÚ��dDO�W��w��b<���>�o���ö�Q1KLXur���ȏS�pǯ�lQ�o��SKU?�&3�1�:�9��}����q$RkLJ�̻��|>ӗ�n�S�ۏM�<�:�z�\��Eo�mG�{s+�5�M�e�R(6G�ՃU��h/k�c�j�cp�*ZEh�	�����I��P����3b~0!(j�N������|en����o�m�|_%C�V��f�E9��"-ˑ�XZW�K��c���	2g�L�9�ɹ���)��f�Ν�?=���+ěӯ��H]3gF�	����[C'�N�,F�����Páz��i�ic�+�2'9��RI �i/w�w��:Y�.3��9������8����5�N�V	�c�
!�#D�d"����搖i�;��?e�xZ��>�˰�#��u��WAu�]]R�Z?Z_���NB�DUf#�[��
���^�n��a4G0�G,F�[�]ŝ���5�q�@:+���ga�Ϲ4��,E$n����l]�(4�R���������I��N�kIlR�@�ߊ����/Mʾ��N0���"��I�Z��S��Mt��y�����h��C��W+�P4Ϋ���9 �8��v��fXdL83K� -ƅ�Ԝw�����)7�&%^�\��kgJ��P�z,���L75�+;��z�ig}��'�R�1H*O�PQvH-C�{t�"D�p`�dZ��+t�b�kDB<���b�0�;�٩c@�7�|G	t�0�e��Ȗ�M���M�Z�WNW�u��[�����e�\���|$�Z���(!��<u8�� �<��̧u�%�(]��9��o��Z5б����	hE:od�F����A�a��(�8���������es
�5�_�oy4��{){��Z�D]3�������AA�d��-W� �c]̥߬5���ُ�%��N�;�b^�6�P�%�����&�&���ITY7���H]z�h���Ý�X��3I��ۣpD6ӛ��XJQ9�&|?��ug�|���F~K6�,Q(j�#�� �h�S�sÒ0��B��|�EH
�-?	9����F|��e\��
�\��m�����dnb�z�pD�9�%���۠�k��D���H�֚�̑C��X�����G	hS��}�2G�^�gf�� ��Yyu�����2��R�C#�Z��!R�L�.��%��,V�3�@Io(FnhN(�jW�K^�%į�m�xO�.��WR����o�?��K}�z�0G���s�T95)���	�s���}W�$#�o6�3��8�$��2�$@2h���*��v5�|�D(���t���+<�"$�u�w��]��Ղ�`�c��!q���Ciּ�n�_�܃\��H�8����F���d���U�q�C���iK�F�=�,�`R�i���.kr�O�deN,(�,{M��K2#��ʄ��2lĀ�b�?gJ����Ě��2k�>�)��;��g�,;�l��I��fQ,,ƣ��t~��iC��c ��kl���-枝9J���#$�ni�����F-+��4S�aJ�ng���@1�DvxA��������օ3Q�}Z�m�_���A������x���'�xi���� ��t��=���9�p���K遲
��cS��4Ƙ���ˋ4�U�:��\�qʜ�'%]]T ��+��IM����@�p��hv�s�AeFH���z�PR�Ӓ��'XW]�֭ɰ`)⻝'��E��}8��{s{tA�H����"k}m���Ŗ�!��e�V8�+��˔�N�e������͐R~��rV��7D��0ck7Ā��+���h�'Q$w�/��Y�6"tX��ɞ�t��]WK�Fg�+�E��u �I�	�y���p��E��٫����� ��f�+�l;��AR�]fy���;����ƛ��_��ub���S��P��K� Oȷñ���?��(��!}*�uj�����l��,sn,C�6�d�$>�;����\?��Ǵ�L;9��r���{��m�:����������5F�eIIr�h���(Q�/��"���3@z�Nǒ;C�uJX���\��;D��%9�i5:hdq�v�O��L�B�������2�c&�N>-��~4jd��1����k@�vq�1N+.��g��W֪�	�=��M$��2-����v �S�J���㌱����8��|;͜�7��P�)jjd��V����Ҧ��o�N���x�`; ��X	@����5��L���&��w.*"�b��>��)���փ"_t��
"��w9��S#ݡ�Z���lμ@r��;�����N.���`�x��j8Gƌ|��c�M`]=�ݘL�b)n
�P7�E��#S\�����+�24`�%�+�i˧��X#q�=���!Fu3v���	kw*yq��v)̫}��"�Br0�����ڻ��ӡ�|�6���)|r��
;���־��������U���߮!�ڹ�=ͱ�v��O��e{�T��������!������T����]�����_�Ugm�+�@߆��љ�����R��c��/M�>�b�=K�I��(�#��J�>P2�ְ~Em�md����c��La�40��v�}��o���_χ3毵VǊUbV�G-��쪞M��>���/�:|�r���_����x��������y,(���]kf����D6�4�A�3�41�^3����� �ҥ�ԍ�3��[@���`�n�TfIq��YJ�g;��\���;bXk��O��3=�L���*�����,)^����-	�P���l�ε��;�ׂA"�a��'�5��Vq&��-N��Z�-X�2WI�B�L��ssSnwG}�y9�=�I>�W����T;���,��O�β�dG}l�G��X��$+��X�ю�~"��ڔ�!�p�j��R糝f\'C#�g�U����M���s�_�>���9��v��a#T���!�I��"}O�'	�xO�`���5��?�_*��t��A,��q�n3��rB��f����z �c��R��pQ೾2 I�5�*K�>
����>�G�:��NŸ���� 3���D��[A<#��K�`����	����uGpʎ�s5f2��T�c��\��qLFyYz_�����Ӱ:�=�I��q\��Iec��Ș�֧�U��z�J�dS�䰅��n.W����tՆ�L.k�螰�H��faFCl��'k�)@C*S+X����Y����#�QO��Mv&U������l}���n^J'���V� �0�c��x��P%+V�o5�K�ϯ�����;n��s=�I*Pȋ[a�d��W�̹��!/�c"�_1| �~�B���3݂�����?��B�xc�|$���#� }�钱p�+����D,́����Y7�$L3
�ԯ���E�"��LR/���遄V��%�	���>�$x��yX} b&7�z�S��T�@^�T����%m���������QL���ͷU�ej֕�Lh�y�mwx� x)�p>y�����+ �E�,qP���Q�,XX�����KS���e�c�1G�`G�\�8�-����/�x;�GI*���ģjCh�^ld�6$U͂��u�=Ġݚ���Ǭ$Po���^" �?�-�[ЎWX����»7�MC4Q�#h��E8��o�'�����*[1o�]�����;4P������ֺwye�aa��8D�`��00I�L;gRW�&g^'h�&��M3k��M~���<���#��|�4�L4'A�Unǫ����a�ɺ�4=��o�(c��3�����
���nN׀e�`��i�8�m���Xc���#]:�3�*d��ƈ�f����P��Z4����(-�^?84��Gcg7���fq=D!�\w��J�|}�1�G��~��b�6\�*�M�F�v�>��\"7eB�}T��X��J$�w�,�?x�(�Ǽ���x��7�G�J������FY��s�&�[����	S�O����rڹ�
�!�y�ܸ��@V~�'ͽh��ʚǢ�oOT�'�H���3����zǛY^��8	#�U��SwS�	���HEh|���^�m������7�*&>;����28K!ݖ�?�
x���h��1M������Y]R���+�@�a~�{"�E|ސ��@�J�d�F�B������p������q`�Y݇<̊6��&���f3%	��\i��Ew�i�]>l�q.Q=�\�m����� ���`����*��+[?݁�����\��3��9�yϲa���]`ڐ��f�R5�*��X�S_�|�G�kݰX�tf(*"H�m�!�Ғ�V.�.{���Dh�� ���w,��F����R�=�UjE����������o�4��O�b?@=�#y��C�P�`��~�*`�"��N�WK��&߽c�Q���׬a� 53�p�s�A�9����^mn���8�XFRs�f~�Gd��s���9������Җ�[��E�ʐN�}��(U (���f��Ҕ[�;J����s��=�X<G�t?VF\�W��3���6����tOp{��ε@U�ȃ��v�M��w�����p�
N�
���v������j����P���2����)���W��mrñ��D��"tH�i�8X1�ߺ(1z>e��$�"��~UU���<KYN��"n��'�w!
Fʵ��)M��X	��Fq�JjGw�s�[7r�GX�Z&A�e�x+v���梸�L	L!وg���hw����<>�/���޴�ȉ���=Vj��䱈�ښјf/E�b<�)z��a2�F+7c����QK��6`���+��=_���F ��?߆��!V¼�ܭ���/Qň��|Xe�'*��&$}����=ݰvhO���T��(�f��zt2���+�9��x%$�V��I����g�I�pǱѻ��e�"���� ����k/+���䏇��Ꙫ�;����<���-�u'2 _x�dE�qԽ�Z��%��`�%���Cd��̟�.4�`��-r�椔�{�^0&���;ٰ(MV��M�̅�h�;u 	[���R�!�G���o�7�O>��q�	����;Lq�-B���,�~'�?HPZ$7(��Me��8a�{CXc[l�1WD��ʁ�E�$d�ser����vǀ����qly�ߥ�'���B�hsA����k�41������J'a�2���4I/����0��9Mi�hdz�7��^I����E8J�-�K�%0�����ջt"�O���4=�-���+�I�{�_NQ�����o����sQ�qLb��2����z���[�7&Ѷ6~��h%��#���\Z�?6�Z��};K��Xp@��; l%'�1�5�����L��aSD@�I��7�Уm+.�� 2������|;�o�$z�檶c<��s�5�s�e�E�G�Z8W��l��"%��}�גV#�KX_p!Mg��9mIA!;P��:ѷ�~��"@�K),kT0�ZR�/��>��-mZ1���e�-�ǡC�>��<���2��-�֚��!X����������p�Ùa�p����l�C�Q%�S��䏤�.D�8���Gn���8�	�˾u�(������B�	��%4�۫���<n~��D�4�Ü�ֈN��`M�#��X['�1s�,�$�+�-[��w+F�}�_�}w%���[r�2�t���y�\��"D5?h�g5b{�j��s���IIQa����
�.\�.9�����Ǉc��5�&v{��GG���H&%�+�tA�	os"��!k�^4�/j�GRKG%�d�"9d�K�R�7���e
��o�V+k<:�L�+��>�?���tQA��-p�-��C?��C4ŷa����)��F_x�h�@���DX�f[����(cɬ�po�'�YZ�.ﭙz�5b2�����O�Pz�@�Ȃ�"�ΗNd�gÃ^�թʨ�خz|D�@�PC�Rc������}:;&��_ȣ� 	)���x��O��#�;M����K&��BV�h�� �-�ir�䮾�5�_::�?J�,)������Vm��\E`��X#Z㮐�Y����}��X恨��0���O�����@l�OK�\�Oi%��f�֯�����:��c��r���[���_�
�\�h�Z�k!%�#�����4e�6��G������c��tj�]�v��:ݶf�T��[V��<z�yђ)��׭UE�z�a3%~ߑkޅ�N���d�*P�}�r�j���j�����C�J���i�7T×�Ɇ�1�@EѸґUta~�8p9�+�z���g5��\m�X[�,!�L.6�CH��{����{�"���o���7��A"���J����ub��Hk�+����Zd�e�Ԡ÷H����v�3�(EP�*����׎�0a���.{jx�Ů�r��[�<�VP�WQ��T�q�1��\� �a���lM.U��9C&j,���m ==��b��S��:A�#�jb3J�P��d�)x���B+j�l����s�v�hQ���U�:?F=f�FR��xO*��"�Vnpn>�!iSc��ܸA���0���+��+����W�4D�+��e�;����� ��ɑ�?K
O1��~y�a�HBd ���d��˴8�
�6�<@翜p��C���UN"���dʹ�Iu�����EIY�aг��('��(`A)�p�ԣ�|��q �K�i��8�w� �	�_��kG{Nv��X�B���>l!Y.<#B|F�l"	;S���<jP��0��q�|���O%���fκ�&\�ݯQ,�Ko�@�ޖ&�a��jG=�c��H��8H0�j������iԜ,7X�׎L���Z4&eY�(R��H%%��e�����2χ���!l������{b�:$O׷�.C{b�<�,���϶�5������׉ɫ�NȂ�C�u�av)�7"=
[���Ů����rk���m�mKWF�[��u*�,�� �.=F�K@�����菽7j�T9������@|�M=����c\�7%�,�%5Ɵ#��dV�R��\*/͎���L���+R|��	Zڴ_����������`��l�j-���5de�i��Y�*��ʖ���T���^g�ڴ�1��^勞�G����G���.-7���� Df}I,�= �9�� ���XY�+��{(�1F׈G�}��r�e�Z��t�Q���/��ӤaZ4
����T��rg���bp ]�^�}�����b��j����䡻H����\%��9��㖸����g���f����qp���뿕T��k���˦
��A(��AV���'?�����"�MC�0�3ПM��w���ćG?�u�`;j���?�ܮ�EmIIX�,.v1�x3-��eKx\��F�K�Q�}�
D0����	�(�A���Fv>O��ҕ�LN�KԂM��sS���aj���r���<S��Ou�l�٘\\Z��9�D��U�6��3�T8躽������2�ƛ���z��6.�An���HA�2q�פ"�o�4÷�����&���":mx�1�$2 �N4a�qS�EQX�FD1<��[�F*���됫v^��(�� � ��F;ݖ���^p0�>�~,g;٠X��R� ��^��� B:ҵ��1QT�Z.�d|�F%�y L�f�n�[;���)��Lg������������N����y�1� 
�Y)9���ε�֡9���ِ�� �4�o��V��a��K��o�c,NMᐆ��ޝ����Eܻ=Vm��:���w3���m�t���Pĭ�F���;���t�l��xj6~�8�y�,�����Os=C$<2��J�������?^x �G��7wY"�������uv�-�[��7¥��<#���C���#:�1&-��q���NǇ��Q^?����THU�����A8���-,��^^���t���i ���`��9��^�C�1�a�Bن����_�s�&�=�kN�f��D����Zy慁d�DL28,x.3��1�w�C�R�ʃ�w��T�~� �]��*��}��T'rσW�8�
V:�:���#�H�>0��'�ȡ�n��J��FP�g���RQ��깈��w+_�ǥ�&n�O�OݚfLܰ�?���;����wy=_:s����tPoƮ�9<߭r��{ y˂�y^J�6�_k�u�-_�w�e��p�ܙ�]4=f�ه�2_�6��B�����K�*�8���[re/ǰ�$\]�@��%K�IԜ�	�����}T��`��
SV׾
P#%^��%�J��8m�7���"���DH�5�O�N�Õ(����7Qnݒ.	�.?w� |a�]+��_T�>�Ċ޻��![w�v�6`�$���C]��ܟ�d2��91@��
���h�0���p�� �8Nd�~�Qr�Q���،����k�T�]�$$G]Eͣ���H��e��o�o�h����	�Qa�WQe�7��濙v]��V�1�#@�]q��(+0*��k�i�n$��J�!��ap:0�Ϟ���[@���姕z�!
3�.13�
�g��f�<u��YZ\�s	MZ��*�T@j=�+ŋ�3t�K���;�`t,��EI�ô�љJ� ��w��q�:�ot��1l��:S��C;��AY�����yV�Pqg8��r٠�����Vh(�@�d��}�>�z\�ՙ"P����G��N���M���~'S��젿�ĪC���IV(���fZ���ek�����қ�1KK��m1�Y��[fQ�A�
�h>���
��u�6�'��w�����y����aTw+�� 0�trV�I�u����9߻y�����)w	ŋ*PFI��ϭ�tw�
ꛉ�g�}"n��a��A�N��]d\��3����ʲ�,D%�P�`@(�b�?v��t
n���9;"��!��N�1�v��0���bp�kA�j8[>u�dsc	^�M'e�⼹̓�a�%;iD݄
��>�|��n����edI�?1Jvu!K[PѦ��M훗��v���8�t��T`����bw�B-NW7�pae�7xhȠ��Lhԙ��[�d�GE�a������䊱0��[l@���u	J)S����x���G^�X��w>����&�����_rXQ����'F��R1E	A!�o¼�.%c}2��L���r97����l��D����0�]}�66H��,�$�� V����Θ�2CSw���YaZ�5&o��Ț4e!�fv����tE�@^g_���G�]&�����GY�p}�*�Ƈ��'t���#���{/�(彤6
�Mm.�_1ë�&��u��$L��}LĈ�M{���/�2�G��#X��Q�V��J�Gp�Ґ�2!��6��K}��;Y������~��r>���3e1yqGحcELq���������4��E�����Y��rJ�.��Q�t;kUV���~�wr�Xc-��*H�pC�窻gq�4ʧ*�з���P�L��_��"��3@��`�P*�"�U��_���*��_�~�Y��SS."s�x��0��c�쥱����Ȑ���K#&5�D��d������m����}�Y���C�صa�k��v�e���&"�+¨�,�^�ER�*q�}" 2�^D�uk)�f�عh@�7�L�,���r�i��-�}�/�±�֍ 	�h�5C��������	P#"R��򩤣!X�I7��SmQ�kvX4�s�|��V��|�	��N<\O!%Д�E�����t��v6�@ؙ���S�X�q��qQؑ%��f!^���G�2�r�eL�B����ƣ��i'���j��}�'AQN'^�}V7U*����s�@���os�N`���j�m�v�!p�0���4�Q���!D���x��_&�Y��$���KP�����$���ֿ���|�v��I�w�<ߣ����RnBO)D0l�1\Y�uKT�����Z�-�4�R��Q�|h#XoE�j-K��2Q?��n�`�	P�C��.���=,6���|�i�nI���-!���Z&�{�����~Dr�W����ӎh�_�<*���m��k� .��SW9с�Xz;����/$�
�ɪ�� �6� L�"�
TqN��>PV�'��S���ǚ�~�����P��7(g-��4Z\!Y�3���~P�����x�X�CĂ���5�3PF�U��U�o�tm4��b��MA8j9�/��8�ki�N���ߪA���|�鍋���P\��7���6]�BZhH��+ �}����VN��c��L�q-���-gzߋ��G��+����,�؇��vo���6��E�G�G����"��_�+��6����]�ϵ�("��1�M#���E��!9��H�]�P��"����t`+�~U�G�6���Q��լ��}{l���G,N����Ս&]hE��)� ۞�*�E�C� q��R�sAw���e+��n�-�"�Ղ_T����nEv~��>�S�*:�']��nb#&�
�$�j�U�mI{K� 	;�����y�AՕ0�!�UWEk�n�KY$���b%�o���
���x�+@BYM�"6���L_~���e�藜D�Ħq�W��'kԤu�����Z�u�_�
x"1���V��K6y�0ɼ�gv��o
�n�y�q�2�u����$e �|�o�I�k�8dőe놐�g܇��R�5�<�,Sj�zX�zA�X!G��Xm����\PD�]Xfm�P�He�&�!tĽF}­&<�&L������_��}L�
�� c�J�= -0������NE'G��d"�X�����h����_�Z���m`Z�A�a�l�ݱP�&X�"��"G| ���k��~�[��Ϯ}j�lB�Q����~���u^d wыE����snU�0 �`���_��6O }n�Rw&�a���ޣfA{� �iwY�a��݅��qz�(Թ��ʱs��~�W��m>�6`{�~��O�<e(3�:�m1,�ӣ@G���X�rhװ�<�Ba߂�5���IZ/}n}����f7��z��<�J��&ˍm�]m�A���L�	�e�
�m�?*�Q6�E/��ϦuUY��<fJ�d���P�����$ ��,���m��w�%����c8���n�Q��b�J���G*;<e'���H�XlxV64EB    6280     f40#F\�Y.sk�1:�<� Me��i뒽��0ӏ�t��Z:�����v�B��~k,;�d��(c.�pI�{����-D�̜�-*����9#S�/�=�ȑ�H��G}*n����_C��8������z���J�!�����\r�_~7��¯�֒ �s,ǎ�&8�e�e��czW��s欧]2�>�����q���ys�k����6�n4�ެ-��b��̒>v��m>ꓗm~�Ba�W`u �|���	����Zp���~�چϽ��l�Ș��"�x����>�N�H��yi�O���G�H`H3���2���^�7΁�y��.�U����{���)Inm�D�tkl�&��_�B�,�w�z&�m��%�Y��^��l��^b��<Ť�E�4Ӡ��uڭ��-�����Tirة����ƺ#H������k��g�J͙�V]��P��hb����n�Gy1�EyO�nd^`ɘ�+��]��U�of�͎�+sɳ��e�c>��`X��ͤ���y�'i�D�{8��
KG?k��Y�eҹ9�����bX |���1�� x L�O�o�LSQ�t7gy,�Q���tB{k��b�е��\�Ty�=2�I�K���̞!�o���|_�{��y��[�Up֋&ƞ��G͘��<�V��w'����vqREH%o0��"#,�I�]��8�p|T�_(_ةg�[�=��:���t��V��8�΢�x���gMc�no�zo'Nr��E\Q���ǅ`/����y���;!���.����J�,˻*U�V�Hߎ��e�)�	��<�'Є�`��*<̃�Bt^����ę	HUHX�+"����3?����.��Iafp)n��.X8�mPKx�?9����}����4U�b��YR8%��k��r��4�c� �N��_eef� ��]^)gU��&{���M{��`(q��������PۓXMMX��mT�F*�/}��G'D�H������c�z[�2�N�eS��򱯝�own���k�D�e;&���ȧ$�Y}9�ݘ���H���"���ν��?w�kE�J7�c	#n����#&�OY����Ij��	�Jdf\Jin��}��	Y�[mY!�GSp:u�L�`2�e�� C,�`I������ӓ[`7�V~[�c���r�*���o�����Э�J6���������g���B�ĺjvr[���_3H��%�O�cW�{"��Uqb���o>��� 	�%i��[D^�Q�'�{h�Y���mP���9����S���?�W��]~��T}ADg�#�4~i6�'c�,;�T88��w���6�aS.�ᾐԊ�y�>3��gלc?|z粥��Y������Ԑ�zs�0)�;Sz�����:u�k��6�!O��/�Q�Ήm	����	�$����7�m���M�KC\�ʵ����n�l_�p@J��m+���a׮��E� pԷ�wK��z�P��r �?�CQ��2��l��	w��h���}_I����[�r����@�U���β!._�5zmջx�qŀu��������J����7@L�$��c\�a-�D���"Ѩ��i���[���R&Of�}��h�[���g�vz���-��J���zS:������Ʊ�aR�c��|��QɈ��%-Cxf֠��:�-���������OhQ�7�m�Bx���x���"�v9�2X���[��0z����[�r��U9��)�����ɥ')�G�鸞�#��ϋ���"���>�bJ����ê���_c����N��N�Z]9�˒�)�T�r��;kr`7�����U��V2�"�b�R����� ^����q!�l�J
�'�p��}���`68i^tx*�u\�_�s�S��c���z�\��E/
4f�/���ā�t���ňC�����j�3���mch�u���e0�7
l���k?����+N�4���&�ȣ�#��e��+��*��m`)r
���a�u}��[%��
�po@)����sD��IbS� ;�g"��H]
�̻�a�&�v�e(��	 ��}bv�V���qQ��++�v6䈠{f��O�� ���v}5X���iPaA�ie�[/+��S5�)&�`$#�E�7��I����o��B &�ו«�b��|�f�\<'��7���ǁ5�v2���m�h޺�j�&d�ݪڰE��(���ʫ�M(,!�4G����fb�ԭJ:8� ������վ�$�����C%*��3����֯�)��%�d�i�ʛ����������p�)\�둪�<r
��bz��Q�����4��\ҷ�	)��m��,�O�M(H�Z�C��θ�L���Qhi�T�K����S�� C-�x"��$�d������e9���%�$����� ��nW���"�U7#��.�*S��D:��@�HbSD�#K}pL�9{�e2j�,ڱ����P��m��ޅ{�v�W�,!y8��cf�R�t��Y���4'T��a�W	x�7p�e���t�8Կ"[bG7k�/7>vm��̼o����t��Z�:w�=�&�u���!_�5�8	۰��Z�CE�ֶ+�F�I��e���W0@~�� �f�~�5g]�f��h S3`�2Y~����9�E�)��hǷ=�ȸ�	M��I"|00�t���>��6fP޼�L�V��}5�[�P:����շ�q�6� �hJ7wyU��&l!�!Jt�%�o��*R0'X�����O��B��o�Y��먠���#��c��B��0�����ս3FR�O5�kͶ��^Oq��O��h>t�;�a��bd��<�U(��q ��uך�֑�_�Ѻ6������P�>_��a^�V��!-����Q�r !bJyM�)/���� �1馪{�,Sn��ȡ&`U��i�ѥ���4�J�_�N"l�"���.�A��[w�ǰ�ưe��y}�%P�j�er��'��Z�6U-o&yp�y�C�R�iPn�@�VE3!)�Z*~�����_��M�j�:=jr����<�-W(��څ*$�v�6;|Hg�gx��܎��IA%t��&(sT���$���^��1�W�
�=]1��geJ�H�A��\��eQ�o<�fp�	L�E�]�։ڦ3F��ea4,�M�����O��,�+�aX؞�"�ҏ�g"��j�(
���5)E4L���o�½��/��zN�扦�P��M;f<-��g��6��D�ۅ��m�W��8��C�=
��
�nW��i�?�pO7uY!H�-Gi�_+�+�$b�	�2?�:��:�U۞d�&)aS�� ٴ��Z����D"6�6$��qEĺr���������i���X���
e��p�z�H��Ͷ��
`�?I��<aWO�/��a�z�Ó�?R���/�%d��ٱpIx�!p��ւ�����c'��6���I �+�8���C�B�ċ��\�ƃ,�O�IT��Zh'x�̃����d�gH1� �Z)�����,""�	��d$ځ�K�6ϓRX��K��t���ca��&��@�GI������|J���?�ӭ�?Qk�>�߾�ëJ�No,���cM�a� ���~͓��?"}bs�l�zvp�ռ������ak&��T��J^�u�BY���d2��5cr'P<���wjN���$��Uv�Nn�l%W�8�t�pD��b�����l�J8���@x� v�z^ge�n�5@����M��Y2+.��Ɖ�T�ٔ�i 4�V�t����c-[q�z�,���ܻ�A�3%?)!<�6���c)�zHk�����0}Û�~�T�V��|�]�?=��P��f���ۼ@m��9�m�q+p��8y�