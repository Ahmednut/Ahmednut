XlxV64EB    9840    20d0saf9����	�������V��%ޘOʽ�L~	G�c��1�[K]��k�I�CEl�
�m�-~!r�Us��HP���JA�9���md�g�Sv=��[K�eȬ��~6K-��hψ0�ʴ8�J�^m�)��~�Ě��7@8�;(/�Y���3㏅{q���r<*!���יM��=�h���P�K^���gE�[Ą����/����_\����S�RZ�h����ܵ���-��j$+�&*��uݩ?�����֧<���ڂ$�)A/&o�-a��?�߆'z����)no�I����!����,�flXeEe�ʡX�=�J l�2����f#`>*ѩ�����i� < i80�2�����ƉW�1^j�Hl6iv
�A{_wVk��]�X�׌�<s�%,��ب�������AZJ�T�SJ#J��*kO����r�}|�`v��ʚ9K����&�����Du��jv��EaA��<;8����Q	X�o��WQ�`�;f��"�����������f8()�H$�m�a�m~gT��S�2�o�2"����`�g�)�g����[��R�|ͷ~neߧX�@��М��6%d�
À0M��S���K��qG�S���BX(���v��z56+oQ�q�&9��0f���P�Yq���}Dxt��xI(+q����X�g�x^݂)�1;.DZ�j\)�� �p��v2��#T>T��t������B�2����bup���,��]#���]L8EjW�b*�s��)���\���vRD�@�|����I�^�m���('��	�ρ�گIh)k��o1��D�Y��-��4�J鬚<	)?(D��8A�������.���+� �*��B��i<y�!lJ�+~d�C����їL
�.��_Bx�V�8��C�����t�܀C�M�1�u�p`�}���1��!pT�-��C��[���S3�1G���T�Y���͌B�����sj
k����2��M�U����!������벽���7���T<����u�O�����y7J�zvÎ��ҽ��(�h1y��D�gdZ;F�ph���0Ł-m�����\�#��N]XM��;��'� �����|�۸�)p�3���GQ�� wߜ��]��2��|J+�j�3a�nB��f��J<!es���D�����wB+�L9���I(5��޼-�����K��2�@�õu�V�,E�в�ܡ��;�be �B��F��jR]]�{a+}�P�.�����#�_���aݛ|�T���J�n���()�1��yU�������G�/��k�2y	��-h%QR����t�:Z�f����qg�ָ��B�W��Q�����kL�x4�#�8���/�7K����um��X��JQ���GNq[�˰��"k$�J�E7%�/�51Iי��&`ކ%Z�i�cR���ک��*0�+O��-����Ὡ��lȦg'����_���d`�����m2����cϱ0��7�
�C`-hWM�mk�Z"m8�+���d|���=Bɻ�G2�Ԅ�^O����l&���{���I:�A��n|6�� MF����Ŷ�Չ_��e:����Be}��l�?��U�{���'k����A7SLѩd/��f�LS:�'p!��;]'Pho*}�uJ��LwlN�`��!0L)����ě�~��x�B<���G�J@vT�0r����D�c�L� ����lm�3�ec��T��۫������j,;Ը *'��2�̂E����՗,N�J0��um(/{G��
Bqw>��a�Nz~Le9P����?5��l"��e�+���C�V^���)E�X�K�)Hd��+ږ�'@Xhҋ&ڊ,���+�����g�����y�	�	��q2H�%+���pSz����V�$�M�����?�Z��-Q����в@�>K:$����@j�d!���Z�nj5��Kb�:�Os�Q-Y�Ӕ��$�rS�pw�uxη;�έ'�oY�}ْ�%��>��IX"�I��z�i��=v��?*4�ç�N�����M�ؽ��,�ѿ��{Y��H ��	�$��CCzo{�51p%��E�L`ڹ>rd��Ak��\_	KLD3��/k�]$0�9u�m#J��8}�Nc�g�u1ڍ�X%M,SG���0�pbp6�)#�,����GH}��:�t�C.ͦ�*��1����VZ���II\��:J����~N0|h,���y#Q�҂��.-EV!��<@�zC:�5,#�L���6��a�64Õ��˶3���)_�'�5�X�������W�������~�G����d�4��qo�i����d#�����GJ��_�>MZO�����"@I�A>y=xJFڏ��G��wS��E��n���@G=���FˑM��i���=�iTb�*%s���,f�����vy-�
lwv8�.�4�:3�s?BaR=l����|9y!R*�� @�l]ʸ^���9��ho3#�qFF#�{U��,2�>ۣ1&���x�REz��]�&.�z8�׍]c��B����ݯ�E�&{K��{�i&���e0.HkKt47Yq�]0i5���Ѷ:���f�x�=f�_�t]z���L�g�D��%���u8��F�%d(�<�����������B�#��a�>��c�-N�i()]P��{�1�W7�T�Z���a��C��
2��fM�P�`xm+S���ٯ�A�ʹ�&�Y���&I��:i���J�r����B�>�;oհ���W|�v@��=,"�Й��cQ�#��1c���d$eO�?��e�z�ۘ�@��V�_���X���&�l�F@M!�;�O����.�5�p%��!����ŭ[�\0�E��~���B�lC�9�9��j[�h�sT%8p�=a�E��p)�>n3�! �u�����s���Wס��<�F�{�W�Ĩ���!�}zs�!�9�qi�F(!��~H���K|�V�]�򣼨ܖ���I�&��{�&&�R�c�r�nk��� ���k8E��4X��!B��2-���BxD6W�5����o����h��n�x��Kn�a!�
����!]��Tq�a��Lb�H����(]�n~�橿�3�*fV}������jVWG�_���7�Oc$F�cf�fA�ˢ�t��`�̼�xv�y�4�sض����Q�a�Di�\ �b���K&L�ݑ�����:�̝8�Ŵ�C?�$8O*H����띹�
,�C�����`��4�ѷ���������Ab�>�e0>6�a� �D�M��<[RUBA5�H�!uX#����nRx.�dEP�����QԎ��05�P��`����A'��� U�z3yu���nz�2���Z�7���Vl��Z%�\0bzO�-9�\4xzg�Z>э�*8j�	E���mN6S����xЍ��b��Ss�0c��1�Tg{�N㽅;R8_���lS��,�6!���T�E�9��*�O�{��판ZQ��ԍ����o!�=��������0H�c���#��
@�������پ��������D���y��]���˶G���0e691J�8r���=Ͻ�^>Cwʱ���m�7,�I���I(��wt�p�����i7*{����t�� Vx�t�I�0^+b	~�H1p�F}]΃2�^������L�YQ���^�dB�I(�H�A�F���\�(��:���;<�h�wϴLa��(�Ќ#�Ot*�T���	Ng!Ȃ͙��԰�mybZ=�u�گ�zX,�.�
_S����+��*�xŢ�Y�>��������$|�t���F b���(d¦�����{��d�,�D���.��c�$C�q:�:�&��㒵�z��&n]m֬�7�#�#[�>���b�V``��0�Y�ߎx&C+#���{�O &��f�U$��wX����b]�62�Q��GJ���ڵ�c~��VVe]�!t�ciL��f��7}���uz�~E�0���*�V����0ڞ^>�B�jj�H5��䚤X�tI\���*ƨ�8�j�3�z����z��TDZ]�-�[��(A���@�'�T�� =o�F8��d��<��1�q"Kb�]��4@���b�B ��Ć�Q�C��ClM��,���Na,��z�Ǥͣ���R�����j���Ѥ�O���!�qi2%�ұ��+�|����]�$f�!-���m�#��y�%k�tX�-��ۨy]1�.<�� �қ��ԧ����j$S��#��n�(�O�7X�mM�&h�H�����e����B�W^��y�G-M��!�}�5���	X)v�%�ʬ-���MSB435�wm؍���N�+�_�Y�8��$��n�^�І:Cj��>_2�n��T��{#��5Ϸԋ�3I۝^}�BkAZ��4����hߏ��y^Uѯ-l�FyĖ8��Y�lXK����Ǒ�#����/��^F�f��{��P@�Rfç�:��*E(�cε�]�U2Zo|��Sǋ�q�HvO[�96�\;���@z�����e�3g��sJCG1��J�������`�T��ҳ�tJ���6T�)>?\o�:iE�nů�s�xh'�]o]��;P�J���Ȍ��z׭B_-.��1����"�qMs!�1)�t��{kAς&�Ѥ�0*r8�U?�qQ_V�}`���;~��j�N;��ҷ	S�R�P�u�:�r�B�C`z<����Q�E�.,"*��F��l���K?�(���:*������H��$Wsy{b�x�(�e��]�}Ph�~���oC&p�@C��$Ј��9t{�3I�'�~ˌ�xB`�|u���F��;`�bKK ���1Ѹ���Tv��'6L`ЈEۚ�� �~��i}��4p������/g7.�d�AևoH���OC9h���C.l�p~�@U��P+b���J��c��m��A�;vӪ����VE�V/���\�fZ�n�fy�G>F�;�ߢ���W�L��
6o�j10��45	�����*�.7�$���{MU���b��-+�;��K4�x�k�vS<x�<��~u��Vc�7�CX�:�W����ѩ�[���������9�A3T���y�G Ť�=�
�Xs��3�������~���}͇�yI�%i�\��!��h�'&�2|,���*�MJ]��X����,0��a�	��UuL�����KI<���?�?f���r�H�̋Ϳ��[J!WY}�<�L�c�%T�������|JEG`��z]F[V��<�)HU����vEDn��L�*_DX����M���3d��Al��U�	�rg oIb�m���<�ؗ�G��ߖB�Q��	\�;��a(ON��z�W}>_1�X���$�"B!<x�&E�k'�C��nBb�����-B	A�\ҜL5��_3>�k!�7G�t��.ݥH=��[f�(��4�i��*�#��[�f/yΟcd�#��j߫y�߅enJ��==����˓4�YQ ��M)/���N3�|5�R+�g�{���Z��Q���Ђ�H>ڭ�Y�������J���.��'ꐐn�����欤<.:@�|�/�*O'�9����9�R�h��[pkc`Lt��O�;�(pPO�S&�qKm"[S��tכ�~>��x7�̎cWK�~:|��<[g�=�١���c'��;-�W�`���M��	��	퓾gPE^�s�lE�!�����?��Jq�>�\S�rHa��w-�#\=�����:]L��#g�{�̫ 3��X\�B���)�A,rV�L+D�9�f��E���X��K �K�CET}��X5S�<�S�[�%��v�5׏��,�ݔ��]j�}!��1���9�R��hR������In�E�;E,%�0������}�rS���Ye����q&ŸA�쿙`qV��W�)a��{[��ǹ��w�}W4�)&3ߊ����p���3 A3����i!���n���fǦHvlw�7��ܷ�ߑ��P�6{TY�j4��bIjz�:_V��4�ʾ�R�~���[�~.a;T�#��ul��`����E��s�쭓�{��i���ì[�5ݽ�<t)��A�r8��q�;��Q��i��R��<��6=�v��f��Å���l��7X�'
#qk��3/o>�����wA{��Ɣ�rH�="���qHCx�V���.0{O$HAp}<U�����opۍ��΁Ҏx��}��@�zl� 6�D�
΍N��ڀMӡ��p�\KMj]�ϧ����8����?��i� j�L�
�.�U�����Ң_ҧG�.<j��}�.��!8�1��;��#�g�bxxE����7o99��hm5�E&B��SH��E|I�,z�v�z\P�3�>�������3�)�o�d�7iw8S_Ki��+���F�kn����8����	�u?�$<Q"��	{�c���U�_J�ho��w�����勤����������6I�4��0G۞�rØ`��tE��ޘ�gm���H����n���s�Sָ�5�P�w�~��dH�Ixɥ���l�q� ��?X��5���S�m*0/p�y����,�T���˴�)�:k��o4Qip���}(�)gQpW_�dn�c���"<�ILFD��&97��&i�fY�Z69*C �sؐ#����->\M�%��:�>V�W���-�{@+��=z3�忱�7g����V���?L�mm<]�`�P�X����I� �u��di��ɓ�9�|�9z)�>�;<Ϸ�HGd�|�C)�϶�2���{v��4h����-|���;�e�^7�Q�V�'����uتӋ��@��k�p�􁖓�<�m��������H��X���,,-݈ �(�O�	ڢо��Jw��7���;Z9��|}�@ׅyQ��W�n��l��(|�e8������EX�/�)Pl�ƴrz33w�]���?��i��n����Y��z�SV'�7cCc�.�7DA]��rf���0���5�e��R�4��d���4������M�_(S	{L�J��Շ]$���/T�ڞ4�0��6���H�=Q!6����B�7����҈�+a�����l�T6G��X��c�ʘ�������`�(�����<�<N���"#N��n����K�v��c�W}Uį2E�����Nؗ��{f2�-:�v�L�z&S/9�X�՘[:�Cs`�d��@�lM��x0U���$+nef%b����m��'�����ѻM�o$�-vW�_�� )|���Ӕ�G����������1��(̻�ݰF�����va�ML�_�u`� �H���T��b�-�6Z�}��":@K�Zi��5	�6�4�/Q��VI!������]��m�����&K���3�huܩ�֙ڋ5=O:�m����rG�]��r���cߎR�3Yub��m��9z�~��2�Rb�JKL@�-�K���1���'Mf�[�gN���O�F�,��.H�Ņ��.Ldd�XXd�6ŀ�,�%\Q�����88�6����3�������U�y?���@���*W�����N|mB�*1��&C!�Mc�0�}-�C�ٌ��Z"�$�X�ñHm�C��;�y �p>��?zgt�54��˥����鬰�=̰�R�ϧ����IT!}I
�˦�����αKິ�N*�zrgɄ}`�#����V��u���#tY�� y����e�P��սX9��O��;�}vf~�|5# ��5���ɳ�3%�'3����nϤ�H���>ƃ�l�ͪkſ��b�3j�
vE<�����ے?K!m
`�'h�ض�A�`'=fݨ��m�h�>E}b�f�����O��M�
j!�_�1�V�1�B�ݻ���N��W��3�z�9��T؎��W:��4��޺�ɘ��ݴ����&� ��QC'����h��^͙Z�k>A}-6ϞJ�n"}cC-��t[r-��d�*��щ0M~�"1M5.����mԛQ ����A��n�/�m�I�w
�FmD�&B$�� =��C�����a��<W��6Cܷ>̞�&���j_1��[�=͚Ν�=�.b�{�e\���?Zh���8g6Wpkq߫���@��^ڥn|��EW5�U4GBqU���m�_�>W�]��(2���ޘ4ٵ!��q�zG�=ϣ�70�=H`t"`���I]hE����p0~_��>k�*Ο�a������>��Y�����g��