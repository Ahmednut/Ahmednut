XlxV64EB    4ce7    14a0�dYk)��:#&/G��D�Np�4WoX��7=6�C9q�{%�ק�?�J�߆軖�.�j�o`�$�0T
�n�n�M���L�3	Y���3W<�U�m�)0-�z�v�`�[du%E�x0��$^p�ƖV�b����Z�D��EӇ�� �5$����+<��I�,�gv�5TGsW���Y*$��󔺶ov��X͸d[!K��4�b��r7��H�f`#1���"�w��1����IѢ�Qr��l̭͞�uVg���W�����R����F�Q�)=#T��:<��J"^?�6����~�}M��T>ƅk!s�-���_������6W2K�7;#��9���W�I�mbZ⭇��CHXPDL���a��,u��$E�(m�ᮅe��C�+"�_�Em��e~@#��&N��PZr�K!6u��Je�2⋕�& �3/v䰱�g�]�_{#H)��Aw���PŌq�l�{6���H#?8�o�v��O��G�m�cX�-�N�*�?r�m�O�03��e`:���R�5x{���%�hN%�C.n2�<O�hː�ʝ5f��~��:}Ow�������	�N�2�Z�I�()�fkL�V=JE����3_�f%�#C�\IQ�$o���)C����;B�ۋ�"[�7��D$�G$2o��O����u��5�%<��f���K�E%��Ṽ�.^�ո�O�@h|�.���<?��4��^8����%�y�a{���{��u�t��y헿�>�������R~��Q���<��\�Z (��Nv�0�B:��.���0��{o8��s�`�82>ǩ��0���Q!$�規�A_����Q����R�mrKʒ��<a�+Q|_���]X|�6dO���;��x�- $���L^y��˘����sK'j� ��жrj� []�r�>�
�w������`y]e;s8�.:��;�%{���&� h�ep�2����d�K�����2e�ͯ�%®�3k�ԅ�҃�7#��ڽ��'��0�BKwpum)}�?F.V,�Vg����E���z���Zw��	�!@���`�
�h\#�"D#k��6[�ň���ܧ��iԟ�g�.dM6�%�=��k�����\��O��ǐ[[��P��)J�ܲ��e�M�?M�I�E��1��]`�f��6+yD���Y�95>�)���G��S�7��-�a�E�f���w��j/�V���p��Ҳ���vA���D�#qk��������im�H��]ְՐct~MI�i���%=I�پ�W�T��(��"�I�?�I�O4��Qn��;ȵ���nic]�1�����@�.�<~�Ī������0ñȪ��'��x*��9?8�����ü���(�z�@�O�N�ݒ_�UӮj����BWo��	`i�N0 �k��Vͮ�f�:\ O'�u��cɝ�cB/��b�y�q�r(�WM�?�#�cRYOK	��*�A�`��v�8��g(��]2�EF@~��,{�jz�1ѧ>~�;�8�T�� [c�bdB��4v�,�=��*�Ϲ����Å붠w�z�	����Jй.�5@�ډ�	�L$\k�h���˼�4��n�ɷ0�i|������	x?^g�}����'��yz�0;)����N;i���ZL�[���u�/�1t1~��q��|M�|	��3�&��$�˛�Ω�ܦ�e 9��g[��v���@���9����c�k2T��+VJ*r�@�b�ͮf�ųe�;=�dS#~D������`8���:�6)teML���P�'�w�?$����������Y��@�{��ľk��P�6���y��k���ٱ�{
*���u��T� �m��q\a4���[{ć"�����Q�>����{�z�SM�'w�9i�]FO3*?w>����#��I�k 0.�������IR����Ƿ�0}F��%綩��)r�������v6�F��x�C6� 䉂��C�c�^`�^Yt��sg���T��ż�X�fy/v(Wϑ�E����������~�v�����dd�;�{�l�u�P��T����G�ٹ<�4~JFV2�I��IC>�d��ۣ��wg+%�w�v��EY;0^�T�z�7��<�N��}F���ldPM%ԃ�����ǉL�ÜD���^�G���d��l��`�u��F?1��d ��j�0�)m�Z	F+�����Bj�:�����LԤ���M�����=�S%��|6'Y�ۃ�et��͙���6\/�i��r�X��9@�Y)�_��6�c�0��d*Ais
3��-�
�b�m����c�ʃl��1fo]��DFG"l_Ӑ��,���M_U7�G�Q�L�æZ�3�ȹH*�?˰Y�ʆ��P�m�5�� N��:h��μ���ea����9w�c,��W��A.9)�k��T�=z0O`���)�A���,���?�N���{�a,�3O��)e�V��ۯ� u�%���1}��R�<� b�a�c��5T�8��o��q��Rf[�Y	�����6r5ry��;6���`%�i����=\��Q�<�<��=���Pzm� bW�IK���=���	N��d�@���l�д|}&X-���!�#Pח�xA�?�m=�:�Do��'3����1�VP잡^u�C��
H��*�S�� >Q�3������	�h���1�w���䅾�~{e��f�躀������F�a~���\��N���|j��bM�d
P�sc�rsi` �aSgLT�z������(B�]�AoS��>3h4��x������
�AV���O�mO�x��dPD�'��дC��߮7��:#r4�#Oh�i�U}8�s��X��U���?z+ŝ��o-G�F�ϳ�  =���:�6'�Fs���]�)��25'���dB�`C��O�7���]=�s�
]]S(�$y�n.�o���C��\� p�J��Н$�˹��r}n@��N�u:��h#��u�#W�22�s+͏1M
�N1'
�Up�fKd@��[��27��y/��<"���/��W�v?�g"�H������}|���[��� vr�-w�W l<#^f�;)U��uň1/���<�O1�R�Y3Q��M!NOg�1}^��X�ĊdnS�
)P�h;{r�g�Jɀm�������-FJUn-�<�m�[�b��>ɌsjC�t.5�B8��H
fh7����q�ԥ� ��|eh��%�dWt��Ջ���^���(`x�/ߐ��!��M0��#7�d�50��6XR���u�A{{��K�ʖ��]K�Y����P�D����\ZΗ8�?��^	��c��J�6OX��(:�߉D��
�[�QG��MQ�_*�F�������:���g�3d;�a>����۾�u�7I� ����S�>�<������&��I�Ʋ���|���Ɯc��:�����@g�WN[fEyD��*:�i���Z'�zd��A:nnqpo��#�c��7��V���Vʝ�V'\��(v����Z9Ң�D�H�A�g�60�3p+@�� �Ww����Ev^�ԋy��6��ރic��?���(s S��I4m}�:څ �((��ƞ�F�<������%�wKJ�"��<���`f����&���F�2����`�C�����(�{�T@���!7T�i`�xr��E�S����텑�D�#�u������Ji�6����U(���|���7"�X4T��.M�l��~'����Z4u�-l�A��=W;|ʆ}>�F����_�q��8X���|p�<�x��.��J�r��Y 9u|� E�hUA�������9�7��N�����=|�*�t��Av�����#��w�k�Νɰ��?h�ZBhz~z��G�JZ�z̛�}���!r��A�҆ϯ@[�f�q������a���c����^ ���<:g�ޚ��!n4��]�C�@Cn0��H&6�5x8��g�)���+K�G�#��. ]�J���X���A�"|z�OB��E�亡�j�Ũl˛*�º׏��39��k���$��/��*�g;��R��)�+�^l��޶���ק��̛pRf;Bϣy���c~g��C`h%X�c�I�d,��>������;9� >����&*՛��MU��q���h��"nFG'�߽�FT�?�h�w,�ڌv���p>�a��b`�54��᏾��N��>jہ.��%ۨ�T������C��K��S�5�4%��E�ɗꑸvx"�p���ğ?ҳ��9��'��s��N���^��j�n�3H����(�]F6V)���1�ȻhS�A<��Q4Љ��D��lVL���ʍCV	�HED��$b(��W�7G�xK�)��S�	]H�ఓyΘ_,^�� ��)���ב��q?�N���1��C������yn���[�0,�U(���	Lo��W<;=��3hw?�`:�$[�%���qcmOV�<����t����OUj�Aɒc�����~_d����G������J���/2s���,A�6�W��d�e�u�m ����$6�J��$�u1rg��^�,��[Z`��87��z�AWYtR\�z_�uxU�E�_�����J|�3H[v����y?�V���]�0�m��C����7��Y��
xǒ��r;d'�k�D��"��᧷��&r���:�<Wt��xr�_̺<�`F�asn�::�Y�2G:�V|�$��)[�^j�l�3�v�����%o�4�,e��h+�Z��RV�.v�K[��h��u�����&�ṫ��������0zd[��v?���$��3++�"��]A�ĳ�b�A�iӱ��g����(��3�Q!����p��&�b8F�:Eh���\H���Ӆr��D:���N�F�ҳD oT�,~�V�;4��3����j�ȈB�^%o��|�zSTz�}5-���~���c��.�w�S�Y�L�{cs��$� 5�0�ʯfx�E��.��!�}i���P ���}��J����L�=�rkW�_5Ã��T��&Q1+�%t��q$����hB�묓��~�
����3����CK,"W��`�x�D�s���Q��v��)��'�;�Yr2Ϙ5ܑr��c���s��('(��\���$j~�b���WuX��>�=�� ԚF
h������!�����EN9��f��>�8r<�R~�y�vg�����i�kk�h