XlxV64EB    4106     dc0oQ�4H�Y��aV��hf���j6֗�����UVQ[B^)��4u�xb��
��ma���аȞCJ��aq��&�TNz=���/����M���6\�P�pы~��*x�`>����Lw�b��!���NF��!�{k������X���$�'����B�B�		e�����j��`��7>W�G��p�%�Z�j�<H[��M��m��d ��V-�4�@����զ��e�&oג�ʉ�Q��. k�yk~˴�gV������mNZt� ����˖KZu����X;OS�-�h�X��g_�5��Z���\w�	�0/�
<'N+X�z�.��l�\�f�+ f[��-�S��(G�f�����2�1-�'��0��+���݉_C�%���u�h�/&~�>㯶�-��w߈���]�W"�f��o�xՓ��A�m9�x��8�Tf\��g���6���+� �p��aH��pkb zv2���I�ۑ�r�~�.���A����+�ڹȵGb��P��OP8|:���<�^,TS���9���:���VZ�U$�������=��2������T(��λT�����5�&$�dgj=ק�L���uQ�D'k�>5��C����[�~�]L���R�?`aH� K�"?�]5P*���Pe�"�԰�<�V�V9���ɊL-vo㸼���Z-Y��{�Aw��f�̙�&�N 1ނ���ʎi��Rx;9��0~mlU+M�&�����@�\�I,���܌.�ƈ��ja���maɬMv�_�3��VJ� �C�$�]���a��:�i�����|�a���ϰ)��` �̿��t�9ޜr	*���'�9�er�m0	6�L���RI$Ck��s���p���hmN�(Ż��-��)H�]Vuk��ʐ���f�'�w�6����li{0��b���*���Z�G2g�B���~�p?��|7+�X&�>�%%bMn%|��P�AV��sH��4�����BUSyQ�~��+��O������!��F)_���`�q�S�)��1�Y�=�]~�
ٶսMḎ_��9�G�>n���7k�_GY��0��
(�y��\�MϏWD�Ӭ��.��� f�3OƜ7�^�$*���iYq�_T`�n�J��s���)k?9K�P-i��ڀ���Yi��Zv��¢t8��)")<�}�+�b�������)�Է�ү�`!�D��L�%��J��(��(�r��V�=d��Ң�.n��B�y�~��i�渣��#���'Ec�B�W��oN��,�i�8l�l���=d��T�@�G��W��%�d���%�iEu*�̂};����h>��%�+�j�AB�m2el$��k��k�g�h�%�Wf�j�ne�6暌4^�,���cC��Wz
�ha1�y!���7�WS�.Иm�J�Y'�iZ�D-�ѬX��P�<R�,���ecSD�>�G�|�U�;�핼��>�8<����WJ!e�>i �R��l���{M=.klkiv��ʮB��lz~ˑ��Z0F#����W��ư=��O_f\�Iu�wVvn��!���_N�_�,�b#����vHGRs�ls���8��:��d�]��Ƙ�peX>��ک���򈯏�n��Lϰ�K�Cm
ڧ���� w��k�7<����xΡ�]˶5,;�`'� K4�?���U��|=�����ʒ�i@O�% =@;�3��n�`o�i�љ��C`T�6���CL^6TN�,_]�m����*۪`�q�@C+�0�j1�)�Ї��yN�Y3�қb�};���s0G�������o����e��G�ʛ�j�Hw��&��y�-幐x�0A���>�J���̄:*y���as�*F#���i�~1xs;�і5��e����k=k�A���| [$%W�[ s�f�7�w���?̀���!v���3?���١����+���\)G��G�?{@�jqH�p!�~|	K�s�h�+�H��y,^�a�=*vc��B��%u����[��|����2�Y_���֪�3����@j���b����x���:m|����vb��,%��!��1�LlJQ'��;M�P΋�/VyJ�4 ���(hI�^l�ĩ�b��D��P���oL�	��9���>PM�,�f7x�0k�+c᱗#W�]lhnu������;�ʌh�^
���+(S���¬wɢ� � @T�k�_�c�PcE����P����먠(�D4�l��*M%�Z�F�E�(Yw	�����Y
���e��!h�`Hv�Ȝ�_m�8��l�>ô�>j#�C�ۗn��R�4tƾ�&��<H��#".K��>�񌐴�:��şt��s�$Ȃ�KnN�G|��Y��c���˷#mdY�V^5�FeW�ď��n{Y�E�6K���0���������,xބ��_��ّ��[�� �lr?��h�txx�S,�ʪ G[Я����j2��'�2N6�PR.�.J��Hs�h�����S����a_���Èϊ��%�}�+^X#�L��G�nM"!F
A����r� ��a��k�k�<����EK�`bpb@ّ������p�;n�Z��f�E;h!�&l�/-�d��Q-~���|0L�OET��H"�����u@ӹM}t��U�Z���'�>�7�;��WQn�Ҍ6:�U��$���Z0]�9햻�����v6����Ϳ��3A�\G�W�A�|e�H!A�F�V�怗��&kw��)2�:g�+�wGx�Yҭ�S�Q�x�����Ҩ5F`1�@"���j�	w�g�J��?�ٹ�exy�J��S��_+|�>ٔ�����Ig@�7y�ެT&@GI�bA�gּ+� C�\��%#v}gCǈۼ�k��N�U�Z�Joe�?�&���`0E���kz�NֺV\�mJ��E�鱧xK����XM�p�;�
b34o�˰���*}������+��82:�7�c����`d�*`��/�m����s bz�����D��9���/��o��Nߙ����:r�r&� �ʚ�"�Ư(���[c��H������;�I��	;I*��D52B��Q��0�/�j�iJ�q����դ�G0�Y�eQ�k!����O_~"�9�,�� �Q��T��@�pOn���`F�u}n�-Xe�_Eˎ$}���]�g��8�ޛqX�^sˍ����T[:8�s��3m�#�Q�t؅��H����Ɖ��A(5�wH�/��ɶ<kE(��e�\��d���OS���v��k П���#;��aF����O9��-���t��U~lZ�O�gv�fц<��&l/�-�m\������d���=�](mH7�Ⱦ�S�1�b�z���{��8�3M�μ97 Ȣ6N{lc��qr?AvJ�����^��-l���]��60LNa5 b��_�xA��(.4H׻#�����׺�t���佗�L������(�c�|-/O7T >2z�J�]��)Ӱ