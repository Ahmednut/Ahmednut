XlxV64EB    631f    1730�9��͠bP:��l��le�cb��<R���e��j���TÔ��q�qr
`^�՘B���_J�E'�i��^���R:��A�*z�%q��/֪�㢑YysJ�3�Sa��-h��α��D�d�kV���W��}N� �Yr�Rw����X�FV���+!���a�z(���%�F�X�TE� P�Z�@��8J�FI6R��#g�潤�� �^T6�s׫��k"�AXA�e�l�]��������I�!�;��:�5?ޠE@$�`˥���f�c���۸2�+���UC��L$R���y��<�k�^Q�r3�\vTݕ��Q?��\5:qKں~6���)_>�{"i��Pyc�u��a�����W��o���D�q�Q͹��ӭ��`�8RNG�[7Zzy$�r	��v*6�ށ}��Q�}�c�k&������JX�����u����|�W"�Hډ�o���-{@v�[��U	��WA����A�J�aI�ݪ������*��[�B�VI�H~oc��@�Ě�i�yGy�v�N�������9��+��	�k�����>PⰀ8��D������<G�ˁ���a����ߞ�򕻥�nC�����
��Um���%�7]b��lˮAd�t�!O���E�)D�̷\ �Q1�R�ko[�S��x|[������!q�Ed��/�7A� v�I��R�̵N������k{���V��s�����7�&����%-֟�5)=�������R��b*�����v���ϭ�;�����BR�%��H�ć�,M�VTݩ��E��me�.%��%\]�H	��Q&���Q�����ڔ�0��E�S�.rZ8�*��n��ԙWm%c��H�%-M�7|n�gڏxq��Uw�z�b��ᕺ5
�>Y�56��*�Y��K����ڗ��nm����+��6Y�!�v�!08�R����bܓ�}� �hxKG�I(��#��,p��3d��37'{;���|I�O��ވ��<�O�A�+m��h�t���@�|�~@G'�u�*OZ��j&87��l(q��ß�S�&��k�W�O��>c]<ٜ-�����`v|٠W��bC��3���و'p�E55�������al���oe��Q����P?�!����<����Ť9�B �ҠT�-AeG�f�z��1r_�7����'�|��۵�2���[;�;�A;e1�(���ǵ����{��4���`����6fsQD $-�����NL�nd�[
�S�R��y���juw�o�`2�r?�:r��)��ˁv�2�w��'xo����Ӓ0Mk�2ޘOc<�?,��2�0i�<�剱���ײ�ы�6k�ٵ����.Vr�xn0_Dn|�*��Ȳ�?��CM�XdyN�%�K�G�i&y1bO��$,�d��R��X��EZ�"\�^��f�H>����5��3��3��uH�A�p��2*z�nT~%��,���I�]q���K�����O�2��U�~�^�
�׹5�h>g�&��&�v���-����f�5�Biy�Q?MVU���q��S��A�n�K����#%����S o@�I,�9�u3wy��+��}�!��5R<�K�cH�^�-4�Y����-.�P��:�r�������}�ԄP��CG�q>R���8I��Rb� :�J�vixC)˟�`K=WZ�����.k5s�aU�� �~�H;��U����x�w��1�Z�����B��9���K�~I{��Ē��Z�I��p/�>���U��F\оr��Ӆ֏��a�U����\P(����y��� � �4+�������B��g�i�����jG�����T�c窒x��}���9M�K-�D�>��Y�E��(1)� jv�{���c�k��a�f nx����R%S��*k�V�ѯE
�{��x���蔞��[��4�_��r3!��	��96/����НjZ$�*e�cx�w>v�+�(F�,��Z���1�,���U;�
�p^�T�j�GFA�,?�n45��O:~�z�s��v���mB�ԪP,O���'��LE���;��K�`��|j�"fOG&�l�<���p�����d��]'H?8Y�Ѯ��#�YOfRS��e;����S��$^�`:*M�Os�M\�e�K�8�H��EI�hr�ƚ�,���+���R�9o�f-"��)��*�c����X�>.����s��:q��P�H�غ�2�?�Q����Q�D��3A]��)}~�)�� �6�=���w�ٲ=�%oXއIr`�.w^H��3�`�y&��A����E-�����D�Q���5vr�`�0@�%�y��狴'T3�8<��@�8oe��M�oܻ�[Ȟ$H�R�л>Y�»E�(;���}����9�K�`��
O�������Ů�5O��L���S�̘г[)ڒ�����нu���5]�l�$kl<�㼓�ܱ�GV��"i�����g� @�3/_�ؿ��S��n�R�a��b�B�m�S�p=�g��,�����\�,JXP��UȪ��U�k�,o�:o���U�rn�D��Z�4�FrJP�%��xi6�&D�8�L{�/=6W��tT�,��7�	>Qio���`9�먕#($�������K���N�0�f�ʗ��7����vR]�ƴ���m��~7�%z�!:T�e���� ��bn�xi�;�����Dn7m^���ł��^X��f �KNB��q�俱j{�F������p��؍�PN�YM��l�l\�	�}�h� j�P�L3�����%��
Fո9\�8xd��	L >!H�j ~�3��Z�2�e�_����(�.� -�^ck��1�-B_����E�*��p��ג/E��%���T���������F�ps�r�Eo����?��_$�C`�����;���!�X��ZW��(Q�i�M���;����+�f8����n\�h^[�)����`���r�:�Ht�ꤽ�5G��<� }�yx��"�<B@E�,��^�����:��j���~̔��a��Tc�<�QϞo��Y����!�#�b�J�]���v��0N� ��qh 끆$�z�f��=cl����x����#BmA,4�W�8����
'$�5��Z;���g���x�T��a���� K}�"���/��@��/�N'�<Ӿ��|�\@��s��q̮,��{���ռC_�lkÆ���Ѩ�Ԡ��Z*�T�b�f�d������m������{��F<R�5ٱZ�11����i�*r�̛@?���`���:�3WЩV�0�0����ۏ�/l_8��VZ�Q�/j�e��H	Y'fJ��
����QG?D��C���:��9eHh<�_T�KxTR_��/]h�.�Wxu��i���X_�J������Z�ztI�A��n�7hȼ7�s��D
����]�c�1X�UO6�w�A�E�	ʃ��.��a] -����[K�8�<�p�Y��Q}���f���m���iR��+a��ƭ��5jN��(JRvg�����#��:��Z(B��L��EH��0e�&��qM���"cU|~�x�<j$'�y���찾5��Xz�di��K� �Ś�]�[�O�OU�I�a���D�G5�q�/YW
��]�m14<�p�ϳp!����DM���{nf_���L=���[�pq)P>�Jk#m3ߙzٛ�O햶�����iԥ&��at�ǖJA�̂{���������m�+������/���U;�<x=�?�ܣ3���Z�`^<�)>��Y�?B�Wvҿu��x�f)ѐ�yA4���y't��a%�x���{ݜ����H����vf&J.�����AP饪�xF�Oe��Y�w�wX7�����x�Nk�x��.Q�8���QB���Sz�������F��}���*B~ռ5��/9p3�bn��3�=��r�jU&��u�}��-Uu��EP��X*���O9ZwS���{��4�Ţ��Z�CCFPNj 8�.�E��%��^P�x5��G�o����4��@�c��5Ev�}F�-�/��2K	_�FZy+:��XT����Tw?@)~pՊ���ltͭ�WN3xv�͓�:��Ë��M��x�	�Ic�GY����I�2?�n&Js��9I�r;M��@ز�߹�_jrG�7)��9��r>p��ef��{�s��m�d��F�b6Fﲋ���O;�"=`T[�|@�@s�ʂ�Ț�}�d�t��RVR�oz(NQ&8/�{�S,X��HT��GN2s�`��1��c|���og�4	���xQ�.�#�^��qꬹ�}���%/HOn]Տ)J�EX�����������'i5O�\5��9�	�ъ�2 Y�\P���!��fPn��3@t�=���K1t%��p��[b�vD���A6���F��k�b+�P�|I	܀5��D"*щ͉q�1�]���.�{+9�&q��X�}0;w�|���~!r �r�K�aU7ddņeS�\�z�XDb��C��Y.����)%�a��p���<���#ͷ*�Q�k��~��%�����8�����\��ԛ�T8�BV)&]��vh��������yo9!���nG&�\zLJ�����w�+G� ��S�G�Ow�)8O��yN��P��׷�.�<dطb�����V{ߒ@�z��`N�Uӑ��)$e.'+�ʑh��VֿY�e(�x��2�+��Q~��>6���0�Uk���ޕZ��"��K���µHW������������*ֲ��zv8r|�V�����zFCͲ�����*V�T$�ͳd�c��� �E�a$�q�%?�U)D�;� n+~dr����W<@y&�gڥw��.?"�)��t�w�����#c��4��F���$`/Q N�G��֟G nW�`��p7	f��"�L��Dd�W��'Jm䲥z��{=��#FU��9�lP�]$��1[��f�˽G]r��ؙ硚}<���/�>�ǥ�m�M�p�:��$�^>�̆��t�N�1�-�+���sb7�G��������[C��A��>��v�#����aa^�~i<��IQs�Q/����UP��QHHg���*��Ȯ��}|~����/����b�`�����G����U���zn��dgE��]�����bi�Ƚ]�Ӷ�>����}������۱C��c7{ds����y2�+o.�*�QG��=�Uj�z����,����x	!��?�V���m��P-WP�Uƪ��g�e�֐e{���Td��:�>�j�GOۘ7Y���+/�8�6��V<�X���3 ��dH�mL�hA�\���Y"�X|�B�X 崩������)�P%�`n!�����1��p�.O�2�I��0V/�g�[���oL�����W�r5�}K�n2���ژ�"�������
�"�Ym:_G	5b��`v��5�4̫�Lk���y�A�����:m�䴔� ��fcHo{Itv�+o}DhI�Ԥ�P-4���;����C�	��w���Pk��5H�:2�5�_��j6s�{g��%��Z�4P�}�i�w���T�����R�34���fL��J�d5��Pe�;B�XѸ	�-PR4�.=��9א��|�"ft�\*�׌Gu�Ŝ�-i��	Z�p[i�kPԮ�t?����w� o[.���nly����ׂ����.����ʡ�b�t��mqEa���e?"��#�����D�Y���T��v%*S���",��Mj�HU�n��sV?"����	��E���h��&�3�ާ�V9t%Zr�ݴ�C���r�|�w�򳢮��<�K�yK�l~���h�X��9���:}�OB/�4�
��>/d�}�m��8�S}