XlxV64EB    588c    1440��御tZè�B���lA�_���d�Zvh�~��ƚ�nH�HM{��I:���*Y|}�l�i������ӓ@[ݑ(�8K����A�i�T�!�ܫ��1�ծK<6sO��ӈ�1* |�*�"�-�`�S3K���Xh=��N)�#��QmĞ��w{�swcȰ�=��}�ר�6�h�)��ú2����	L=.�E�fv���lU8�#�Vb��,<���7�
�rn�5UŜ��׫ز$@��7�Vp��g4�2�e���^���!j�FP�E%t\�V8[d���m*s��2E�N�7��|f��i$��d��/��)�ƅ�,@"���Q.<5��< B�F�b٠S>�cH��A��Sn��Z ��yK��z�h��8�\�#��I������-sw�^�"~`E�)�6���ݟ�&-�|�����D�$� E�����Z��2�]w�[3
�*�C��a��q���ukQzl��c�QͶ���Д��yo��W��Lw�b:��Iw`���8�K┴%��C�;�j���H�-M�{s5-O��4Mߍ^�MrȤ���H���M�Z
|Wg|�*w%��c��vX��arXB��ۃv����b��`FI�ǢrSj����ȌK|Kq���N}�>���9��������z���[p��ിUEF���[�Nw�Ĕ�hW����T�sw�fX�Td�Iy�[�\/�H˵�K��upm�Zd/eC�cv�������`�,�<{�KP�OҖ�m�|9�����$z��q�V��Î��V��T���tI�z{�:��G�]�!�V��}`Z�B���\��u
�h����^f��~/���E>��ߋEb�i�z�!���Q"@~�/S�n�=�$J�*q�]o��w憘�%>�L��W] E����QҸ^���gĮw<o���c2�7Ha@8�3���j���~�7����5&�(�7�9��@���N�(�����-m�ׂ��x�*�`a���pl[����h�0����S��.6hD>�u�6�U��jG����5��s��!X�;(��#�D���2��k�9�#���G:^���cß����;�Rm�� B)0Ƙ��o�xvw�f���,���#�M�I�KHah[<��,��i��	��X:1� ��'��y���<՗P ](VC�sy��P��D���V�j�
6v�zA���ݑ���r�Jp�6s%�!��k��
�l4���UA��Y�s=sc`]5�����A��,�/�r7�ȓ�7�l�:�������'Osx�� �CJ7�e��y9X�Εn��3�[���+�c����A�F�[.!�F�\�~Ccyه+nr#��F�_�c����~�0ŧ�0;���<s���Hf��GP���V 㮋-����J2�3�L��tI�>5��7���@/OHL���f�5C����ÊGtS�\�ݾ��*�e��9l�p��Sŵ:���й!sɷ���9$&�z��ވ�U���!��G?�ϧ-�^�	���M��x��J�	��	*�g<y(Q6�T�ʃ�)U������#�����J��>)�����5�����k��W�-��Dv�i����TH���$��1��%�>}f2����d�/D~�|���d{�7����2��,:���1����mt%U�s��������V:��*�Xw&>�҆d�K1T�P�I"(�Q�T�h�f�d�4���������>�6��!��9�"�MQ2).�;-��D4�;����,��;c�N�e��d�U8�
����_�a�5�Ǹpb:���d;�i��]U�014��`�[-2�)C�"2_$�&JрO0_�)ʝ��e�T�2P'а�G\*K҃�(��K�^�S� Ҋ����!r���hT~�!��/Ne�S��ۧo��Ь�l�f]=B��q�`�Gu���A�W������?I��륇�B3�8ϝ���X�5{ͣC�Q4���byH1�࿘^�h�I��F9�--RN��L���P�� �� T�<����q4XV�6�O���ɳ�ˁp��h�l�M�BV����B}�ƒ~�d�}p����
�NI�[=,��Aa2���H�~�G��lZͲ�N8�
��%������|�eT�}e��(Y���If[�������ʟO�����?��8�[�vIU����$yԩ�hJ��p����uH����n�},�p������6����"�Dc�y}x��t�y�A
���-W#�.M�4��c Յ��$$eŕ0����K'�y"a[j�=-���nS�o��ⅸ{�T��P�V:+��3�)�c{{v�o>Vh���=X�F?T��]K<=E�h� ��K-���f	U���ٶ�-�Wt�O���R�⺲�8ɠ��RW�]�c��\8�̜���Ն���X(^�v0[f�Ѫ�� @v ��5��5��!�[8q�lU�H���/�M�Dx��u< ��x�������u��3"8��-�Q����A��<�)h�g�������?�Lb�[�d�p�(��fZ�<D��"�N[�,���Zݸ����a���hP��8T�����'��Dڴ��"-�yM��9�����C^���Tu�j)�^�� �������O��=�:0�&��Aƅ��{�:���Ro�3��DėKei2)Y1��ɬ�=�Q뒥Sd�nT~qm��l	\<�����7B�ń��RE�9�-��3BV�9�UŽ��n��w ����l���#�Sj]�Z>��G�_���m=���x��*,@|���v?�Ax���Y���l��
�YQ�L_aV*��Hr��#�E�0�s��K�]Ӄk]=��w0� H��.XQ�\[9���d��i����ϭ:��H��|;�שeu1��"���7#)<���BI�mj��r?ޫ���:�0�X�5���MB���Q�A5�l�T�ocu��K7_�x����>����5��r���F_��XN��7��ug�:���y�/]��������j+:�S�Be��+��rf\ʙ��˶B�c�䣠���S���YW�G���p}�R=�+F i�ue`��3c'���&R�?X
��(���:� �e/���yʄ~�N"�/� �-RB�lp4k e�� qj�S�=aP�Tb���kƞu����,��T~��~�謁��#4"�	�z��٧3��e�-j�ĺ_��q}d�N�q�`7<�܌��Y�ʣ§g�h�����0����g��+q���ݣxh�5�O����y�9�s�Q�,��#��EӟP���!c�t�`
R1 ?������X��&��&�4"��y���QAu�\�S2��b�{Cd���\fp����!F$��~�PgO̎�a�p�!}}��Q�/���
��<��4��f����ޟG/��|aH=@��U��ϑ�э_����Q�.�>}/���˝(�K	�[�3gAh�.�+u�Z#�o����⏶�C08Uo;a�/�E*9�߄��,5�K�4�3���.n���f2�صi��#�l���o�!f
ӲG\�g��j0Ɨ�&F�/39��@���#>���V���������JQ��]���_}D�Dr���%�(�h����z.��V�M��-���ƒ����VW��fU����=���*s�!X/H��F&)��ya�z�qx�=AFuF'#�gLoC��2��hd�������ϻ(4��t�Ϲ�n���q��g�6��c	��3�����
�J��u���!��ڛKg2Ow��f�"�-��֗�&]yID�j_d`��59��~>�@�@d��:�<���$اl�BAS�%��M�fC�1X#�Z��ۣ ����We��vI.�J�v��ɮ���A�}?J&K0!!*y�����{Uv����޽�~��pU�@��b��_B���(�@=�I�ω��8'�*UɊP -��<TE)d�a��f-=Z�A�^a7�xT��t�k�Y�e\�s�a�!�1�2	�~�ՙJ����6a =^۵	��P�R99����Б���~�����*dj/�)kjmz)��F��)f�%Mګ*j�]̆Մ���|%N���Q�.� �?^���N-)�4 ��rT"�3oe�U�&��@��`�X��k��Bڄ�w��ƞ>`��
��ز�%&=���rO�أ�����0Z����n1�*���@�P��h�;��@㸱X�3M�q��3�����%��V���1�:
�S����^����td��F�v�HTC�q;D����&_�6�es�)�:���^uFU�����;Z~��L����g�����r�D"����L�#"�3��Ƞ��`���Ǎ/.ϰ��%��8� �ِ0���3��`��3�FK�@���O��g�����������ى[�r3U�QՕ ����An����\�~R&jE��8�m�P�#%�~�[�1���yq�S\�o!��0�� ��p��w<�O4�����Ѫ��ѩ�L��UG?���fj�d�^.�$Ј4�H����wM.bN*#m�^E�aH#ا��گ�-�V k\y��;+[%��<uJbx��՗��q�L?:�^+��|�z��&�s'A�x��K��ݜB�䵨3��C���U5�3kϩ�]�u���� �H����|���1S�!ɷ���̙�nu�����3����[��y��-H�N���㷻��	*u��R��9�T-r�{|q�Ɛ$mb;����턍��p�mM����,H_ގ�������@I(���!�uo�u.�q�3K��#�dM������&�[n��yW��A�P˄����`���U�>����=|Ԧ�:g�a��1l"���m�8����;魼=�0m(��������
�;�����K.��L�6䍯�k�|b V-x^J�}�������r��t Tƃ�U�z,�V�}���,.3Ͽ�K��G���s��<��fh5|�=Α����K�}%�c�i���Ov ��5_j�&FX��R5o�b��5 ����UZ�gM.{'P�Q�	@��I���o�X@�`nk6���DNsZ�l������2��E>�#��L��f���$���K�����c�lʂ�Z8s�1B��h®"�
��