XlxV64EB    8235    1470�on]���fjL_�&�����VP�{�#��q��]R��l�B�Cn�ڹbFw)�b�����C~��f;�k5B�H�ʀfc�K�F�m�)�a�ѧK�A]?�R�7��Y��H�SW^n��|��
����<ݓkkݾ�u��6��T�Z��~�|��`���)���`F�!��rR-��|���t�hz7ɭ�3�^ꬓ�weԇYj�y��ͨu�^��%ѝr	��.�Q!�ASw��>ʕퟌ�=�$z���2F�p����䜙[xA�9 -P�4�׍h�[�:?��mR'���n��F]#sO��זKr��]y��.L�@�����������1�T��c2^+�����°S(_ůH�T�B[��h �Y�YC �=�P(�����-�2��g�������Vo��턀`j(��������f	?<���P��oĠ�N�{� ����a�W7E�?�*�.3j~�?�4V�Tqލr$��H��`����L��X�G��]X���jf����r�f�X3��q�|��,�4U%�x�������8��(�S�@m���id����Fz�����fPJ�q�j��6	�����pZ���*��m,ʏ ��KՉ1&
�E���O(R�1�U�lǫ>���TȓQ��=���b�@1�"�Y�j��C�VZmQ�*
�����cW{�����v첡�:��1��g}��n>���]������G�zK��A�c����[*pn��R��������$��Uj�f��?��t�����m��� ���`8���p��]�71����ٿeDi�uy�R3�߼J�8�(��x������Vi;��D��]�K�}�Bn,/=��x?��1�0e#�ͣ�����$
�2��FvHG�#�Q9���]��n�����;H��nC��ɽM�r���rrN����q�ѝ-����EȭDQR*I�} _�Xo
�g�9�������.�P�N���0 7D��<�O=��X���^�ܺNθ�҆fO�\�b¨s=�~og$�@�eH%�ɱ�4C
�ō�	�x�"A�Le��CO7�H�y�^��w�n@,β �_z��p��K���-F�����.��FS�&�׭���+/6��|h��<u�L�B��l�n�ҠU1{l*h��K1x���K�H�+��b�Ӵ'��2}��x���A�'� P�d@��/Fu?sh�p��t�!䂟1�]rz.��@뢧��$3x�.̟N�W��}��3�{= ?�Wmy7���LUq��)N�S]+q�����ҍ
�����s�^rz���8�N�b��e[ːp[�����u�s;<�����>c�$DDX��9"kb��F:H�I(����AL2�܈L*�amCd��1{����ā����'%,g��HS�i��2�E�H����)��"eU�ud��|W�n+����R��W�����nU�խ]��ƥ�*��*.����ʁ�޼+�vZ����~��ꏶ-�Ot`�}�M)k1�cp��\�R��9P.!����p�o��QL�3���`�t-�ǽW��#ĶV4.��2�������-'I>��ʲz�QgbE�5D!���='Ͽ,���b�h�mzEo��Y�,���~[v8aɸ�oC����[d�6�BC?�{Y��uh^N�������z�W7*���,�ä�W�F���e�Hߙ�6��pXV �~����=؎[�K��h�8�ط�4��*�ò^<t5����A���������\��kjw/� �ތ_+Y!vq2˿��cmg9��h�ec��U�q,�7�A<N1Y�!�s���w��%��H�
	C9�2n�Vg�ip1��U���[�T���`=�َ�[1���E�,>pSh����f�F "�9w�7�V���?W�XM�9�F#������pD�N��^V�t՘p֫���� H��x�G��P=0N�{D\�X蟙��Z$;�ݥ�������W7G��1��]MGFH��Zn�;@L�?]�I&�v^3˫�rq?�`����DG��,̩B�%�Ti0�~��FWl����������ow�ꡱ��J���֌���9|�W]��������)�X�Jpۚ>3�}1����.��kW��c�FU��Y`)��+�Cĵ
���.(?��62tK��w�E�mІd�f�W:�b�R
{�]$͇TQ��D�~��~P+5W;�A(N�	�*���?k�a)�1�PZ�t�B(s5��}t�&�h3��K�Y�f1��D����x!eJѿ�U;�39	(�,p���$�00g����}��z�w��I\�V)ֱ����=~����/WU�[����cD���dk�o8���*�GB�:ӡ����/}#P/��v�«{�$l}�^�lX����2x�����$Z x�8SN�i��v��H��W2���sV��#)�E���	c��@�h썑O��drr��d�mG=?а�!��1'[�rR�a?��f����we	���ﴙa-����ΛJx�2�nө�-��KO��5u;3J��]��j鍲���7ej��-�P@Σ�׋-I���T%>��}1@�e�	�J!�Bk'c썟Tl������,�<=�v�@�Hٲ�.����m��R�RDp�G%I��~�a�L��l|~m�Q+E4��B�>��X���k}}nՒ�.3=󨞈uā
�"./���c��x��65�[Ƙ�{"��~����W(rk��[B���g�@�+�f|�5��Y�Ƒ���4��9(/`�����7���NU�兘�6�N�*�ќ]��d��r��㈺ψ����a�n��}h62ǌ���l.OAѦٶ��'�6�(�dv[3w3�@cCs�k|�c�8�u� |/{�Q����o1�ro�=NQu�������9�k���x��m�� H��P�AFqȆ-o�[ϼ^	}��H0�F؁���f��O�`����dW���V�[���)ua�>�����}���bL"L N�ۑ���p�hcmw�v�,�:ӵ�����EwIΟ����Z��t�*E����S�ML"�C�<'u�~VZ�R:=�ߑ[<�[��L�qV?Q�ltX��y��G}���Ώ�A�RF"t��$n�/�CY!�n��� �Z����]u7.�����k�����#y	���\@">7�ʼ?�M��ܯ�=����	X��0!HcD�[��V˹�Ai��q�I��X��:�WB##B����V�ޓ��Z~�&�7�gRц)�˳�dg=ֶ`}$��!��D� �6ڮ�AD�d+���������ȁ#)�y<��g�r(�9f{'m_4d3w�~~V��|��X��A�/�E�eݚ�i��Qݦ����Y^$���~v4}eQ'pzJ,�F���s�m����	)�b���M%���C��&��tw�U��LE�3�p�%܍��X<���5ѡ�Ԥ��g�"9�(���!T��r#g�9��f)X6<��届�Q��j�b�$�fc�;k�\�X#�* D�%�xa�*�)%���}&���z�!Ѕگ��NLPX�d&K?t�����4G�'���7ӫO�B�|�6es��H��=y�ݲ�rl���5c�-5볠V��Ta��,���*Ť�;4H�u�+�1b�_�:S��y��(%��6Q��$�x|��w�A����K�\�W�P/|��n�J2?:(�`\�s�hI��#X04����{`�'u�/E}���
�o���ﲏ��2�]���Q���9�N8<_���%r�FH� ������Z�6��'c]%�(Z��y^���9Km5re	}�ǯ��K�&����Ѩ�&T�oi���u��S?u�b��r]VsDѷk�*)��������h�U7<��%$):����x��EjQ�s?&�lH�~3m���en��&Y]-7T�H�-�s*�訕�G2�b��M�S	ھ�0�R����K�^��� �ν���1}�K
§�-Q�w白K���)1�`����-Y�_�J���4�A�*T�<��^�.UJEE�oqjiUaԜK�n{�H��6ZG���m�[;7���v�rm������An�|15�,s�k<]��b�Tt��O���[mc�D)�����|�m�����֢eB�����5���	�~��WfΧ>���/�*�KR.����h�[��Ҥ�x�O���"��<�93i�ܵ6%��"�lG޹ڼe-M3@�c<nU��$7��^�qU���6:@��%$��vQ��s-��b���x#%,b�x�Z�O�tcTm��Π�<X.�&A� ��f��@�֜S�Wj��|�%sn�]��Ud�����U��&��s���.��$"�����x�u��Q��jE��"#
��R	��e�I�FV��/�gݼ@ ��@�K�b��������^$f�>^��n_������>��V�����|�������hƄ/�ݚQmS�� �Ƚ�����Y#��ՙ�����=��(�E䍲r�d����`*3��n���w�\�.��붟i`(�KǳZB������*⛉�K��h�ȩ��6[2V���_,L�yZ�!\��P�t Y:�(A��N"�?m�]�S�ӫ����4q���3󯔶#�6w ��a�4��� Q'��AW@��*^��/���o����&@�*t.�-�"� ���8��fũ����c��g��,����䆣�Q���|q���N��W�f3� [R��y�t�DQ�Y,+����q�ڄԙM݋6����ThX) �F�*�:�Ve ��c? �.w���ـ�b��r��>ŀ{\D�f�S����z���.��&�h]8Ioo�`l������F}~���"�	��_G��3Z��5N��ˊ��û�N����?a�����>�\`���0��p���-���js4F!��#bYZai���S[ns�4���j{H���]�w���.���R��)�>OלUə�Dk�S+g ��������5���2�O=>	��c���u1T؅�����Ϥ������_�t��?���@.�A[X��Tew�K��� �9�׬%��;���NGm�m�0�{���uE ��V�����>�~1��yV5@�
�-�(U��9���M3Z��7�yU�c3