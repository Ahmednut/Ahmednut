XlxV64EB    45f2    1160���E<�u(�uꅀ9[n�2�&谿7��+����K���^/t�$�X{��g�a��O��_���i���5�G��po���b\����Oȗa�O$d��KJ:���5����|UD���������-��\���P�t�a/�)��w�d���QO�q�4m�	R�����ڱ/O������@r�8�c�<Ul�Q{XH��q��%b�������IC�a<'W�QhD�c��t�64�yd�r�r��!�,5����������W#�F��ZZ�<X���=��}Z�r��ӆ�o�4�[�U̬egXzߥ�zb��*��m�4�!vA�4%�{X�����3�����Q�\�?מ��u��7׍gMD2)t�=���-����-��.U�=�2?}�#'�NyË��HQ�4�I=�)ZL��NM(a򂲃��}��� ,khd�ucM%wV�*1��>�빛�Y�k��bk�P���Lǐ�8��%�La������S�Yґ�fI�Z#��r~�?^Z�:;F~,U�.�&�6F\�Qs�<_��+7�����#�Ygo%���	�^�eW@�b�
�̘�`i�/S{�Lc��z0p?K������lK&oDE�-�n�����{ki�<��X=zd���<��d+�<q���eGu�Ygڦ�
�'�!�)!>�j��M7���*#�� ���w�� �~*:i0��y- =4��2�f����L�-����C)��霖���T������*A�AAa�ʥ}������M2q"؁5���άtWrv�P��>���WlgN���;���������Z�
�׮��V?���b�*]"S@��u�\�s���V��}-s�!zڐ^����� �&�Z�+QN�~գn��@�o��v��p�ƀ�f��&�;��+�_S%�(��!:B�W���'�6��QK�8u��³���J��݁0x�ϔ��]�f?.>k���_�"��T�yzD߭���o"�����=���2�1V$5w��ԍ.GpR�q�c��^*��G��:�j�4�}U��^��T7��֟]@�R�7m&�R�]��5��� l�/�@¦���mlO�l�@a>w;۔���}�4�%~L���u��"�����xyL���*Y�!����Xm��Z|�8\��	ˍg�[�/��V�ޡL{/}��b/&�\�iT�'���+�Mf������C ��mD��1;Y�Mr�"P�Y%�����z��#���n������0m�!s�(�i�K�lץ^x��S
�h�C_��&B��f�N��d �X��{��G�����[T�-�F��������Hs��0h�U���F����))�S������ti;��3 5�z>�L��w�����Bٴ����G��v��%�g�o�����_�Rl�+�I�^[���=xc�����������S�$F�_y�����)(C�Xߥ6*B�?޻`���^Oq3�7��@���$]ч&�
&ޙiz��ݒ�xt號����nl��w���v%�2Q Y��A0�WhT����O]hP����<��&�"���~��<le�ݷ�%a?��䱥���(�BÄ2�c:?�c/�b���K��x	��]��-b���"N`�*TCr1j�^L+�TaQw$/���N4��ܤk#{2Y��(L�K�׸�^=4�x��90�t��5:�!s}�cG��q�K}�4'Aɱ2�s��7?�蟽�� ��m=�� fr�"i�-sh�M����._�Z
M^#���әΆ��7N�/P�oh�Xmf��=3~��� Z-�R5����|�atW���q������5�tա1 ��O�	z90�����Q�jЃ1�}��J�u��ә����&�H�fb�|�F��M��,(C}����܄��)0�ʾ§��w�ˑ�ɿ�R���JT�n�Pm�tУr����r�[
�M	�[}B4�z�jVz!U�]o��������,CU�wS�Cf�>��YDaql��{�����WSO�]/�z�IM?��z��%>�|�^8%�#=p�%g��<�:-�U*v�D�~����(�#E��Zی®�(���P�,D�ƛ�>��yiнMS��4h�I�� iKe��YZ���c~͘��V\ܤ�҃��ĺ�8��132��xR����t6��(
S窙�jI���Ģ�~v��*G�*_�y��EQ�l�}AҠX���6�|�	���䂏P���F(@�U���%5�L��ho�̽�����/���Wo��Q~(���f����&�A@�sV��;��/��^��щ��Y!��\��Kq��-�iC)�-%�q}��OE�{p��u@r�ąR⥤������=�{��+�.� Z��A�n�����$�����{�U�lk%�6�&-�K�69]%�ܓ� ��ڽM��u�2��.qs�,�!3��N�EeI�Cմ'Aյ�X�T'c$��{jTR�2��a ��UI�?�5gi,|^1�n�����_M�4'��?MOr:�����Y�	�48H��P#���� ����͹)a��m�$-F%��3�}4�,�_�d�޴�bs
��~�H�㉄:��� ����zg�CM�44��~�����L���Ѵλwf����C=Té^�R(�I��x�B�t!��F1Z�+�AV�ax=�|ONJ�6ό-�3/4�"��4ܨ�-��I$�c�S�e��K��k��8��ķ�;�3���i�\H��#}u[�_쌊��kٹE��\�����I�����x�6�6d��j�7N�JX`ͤ;������+
�g��5Z<kʁ5��(4g)^���u_/D�s o�-/ �R��&h҈%�� �H1&������ە+r�O��'�o�5\;�נ�"ɳ5��8��o���k�s�������5�	Jw�����A"$�* ���w_���\�+���L���jaZ�h�T�>��s��C�e����ώq��vG#��<Q3u�r)�҃:xgN�H��q�q�Uk�.��\_���P��]���fH��K�����9�'�	�u9N�e#l��S�C�1?H�`m?�n���=��G�0���_�˳�MEH����S�3�h?g�]s�8O8��Z���Ohy���.o���*��~�\ I\�ʹ���@)[i�F#���u�YR�(WW�� �e�x:n��cO11�N!�����b}~��Qf�  �p�2TQ�>��XD�[�״��'�-��SՅ��!:wF֨�,�v$��#sF;�;��U�
BH�z�rK$AN�âVמ�ǅ0�ɏ;�T�KG3`{��#�~�l��C�<�0�u�:�@��2���?,�N�Ʒx��{��A2=]�1ݡ�-��~+�y��$�{;e��T��p18�1�j��4^��n�k����|}���g�>ls����vܩ;���H���L;���� 㧃V��KQE�i�ӟ�[s{1f��CzJ�Dx �IY����r���84�J�=�&��!)���Xq�WWw]
�u0B�%Q�ŗk��[���0��g�	9�	��<.����`B���.�cɖ]mo#��a���2�Ϡ.�U�������$�6�����U7�?�k�~��|�@�m�ٸ�A�}h��S��F����Ӿ|��~��L˅��8�U�`G��ͦ�Q����/�pLBZ�	�B�4a�z��R�ƌ��'h݁Yl��1�<��uq�K~�k=���ki}��m�q�Uł7��x�i����2ҙ�΄�#D�7����-�nr*Z]�U�-}m��?�� `�WC唤[V��~�02�Y�jeW�j��Wvx�z<EN&jK�c� �fEw���������-0�F��/�}ղ)Ɓ\��~�5y�>��L�k�[�����h���� kI4z򱝗W�����i� -�ޞ
��|D��[6Z�NE!�߾
T���&� !�õ�L��L�
�b2�{?߳�1�,����
�U�!�z>��q���ގb��p�B)����Y��{̺@0=�͛M�.z�V$|3��d�+�Z�Y��nR��tRTL2:ޤ������cؠa�-_t�i�2xb~����H���7�wt��o�$~��d�$و�歄&�c;V�P�v`��^^U@�m_��v����6�[�d��DZ!�-9\u`� ��zv
U
~�[�B�<��R**Q@���R/T��Ut��v�RB�x�rE&�sA�daI�oc6RY��ޛ��M~G1��5�Y����4fi�YF��2m��"���z5}��M�O�� ���P�|�Uh���T	���~�!#���,쿴�ƍpoS��)yt((�>&�M���=��vߴ�Z�	ե��*��x��ra�C
4��B��8a�ڝ�e�A���5���E��fߗ���L��]]�)�����Wӌ���