XlxV64EB    183c     870
sw)��-/8���m������c$���
�f���]��8�蓿�+ǘ{+joZ6���t&ޕ7���&5
.d�9wJ�+o��=�ťHy�߄�ޒ(��&h>������y���������I�1N;3@��I.k��3gq��g<����'�N6���7��J�?͓����T���]��e"����\8�eS��Q�ٴM��x4b��`b�ѥ��E�r�ZyF����9f
`�iA �1Ճ,+�ř)�v�vi��]�Q%�R������i4'�F�G"XR(�fe���'$��3F�g���m,0�MK?	B�u� ��\�όR���{x���XO9�{��&�Aٳ��Z�������W(9�
J�kI��n(6v�Hi��!omXA�W���$�%�q��?F��<)��u-��,y�
y@�w���PRK:]��Tɔ�hY�Rζȴ��t��q-���\&�b�%:�^�u�g��ZNl��K�*���7`�.ߵ��U�*}�,����.�����Es�<7���WI����LU-F �5�]Ć5-�ig��=�����3�*$���,�������h� ��X�l:7�x�"��CyU�ʛj�j1�?E�K������R;C�S�O�n9��E�{;���[1%�+�s �T&�Ǹ��=��YÕ�[�@�{(h�n1�`��]=F�vYUǡ�.�5kqK��3ۜ��~�	�(��Y���?�2����DÚ�]*�՟,�T s�>a\ڻ�H[��GbfmkNR\�~����A-_@T�7����<i��E���@xQ)�m������B)ł֍��栂�Rim�Mw�	�Q��_\ڱ�q`8�v�Ӽ����-�2�_�"Aދ��%��C��΍���)b$�1���Ǜ���N18Ӊ�D���$���լ�ag�rU@���6�,n�榿e3�a��~�g�������h����T@R�(��(}��+pC#�����m���W�� �����r��Eh`�vA�˛6���y���� ���h����,�g�0~>��Au��E�7�,J; � �PU6؎X0!�܄����&�#�N�D�(t�i5��Wvθsb������1���-��o��w8L=2AT�>lQ�
�����塚0��g~�K�W�x��Eu�G��0W�0������ �6�Y	�$|X�����HE]J���
Ǩ�S"P��u���6Ȯ����?�I>���~��aR�7�Gq0�9|?}i6�13���I[y��kF,7�4*�`%�n�n�P�@
�`(a%R�"9cfS{������\���2��j�IQ�hڴ\�KJ��lZ \/A��r0Y��(�i��\�Ȼ/I�=ܰN�ymy�$���g�$H��H=��O=�1����$��K�D
K��qB�k�K��`�-*Yڦ��<�5Z�x�zh���=upJn�x1w\�zS�d��!H�O��"��j̺P�:�XNU��He��;��}�"C���E��Y��Qt?��<�L��[�-ǟd7������b\�0a��e���R�w��ۣR�f�a�B����-��W�O��5y�y��ȓr�Qo��,W=/�x"�;~�>��{��<�3�}�*S���V���O�>5���!���_L�~����r��+�5��yA��nZ�5��l8Ѵ�� \�p�kTS]D�a\���E�g*��ס�:'�'m]\Ӿ�~9�2^��0�+lQфZ�XS�Ww_��z��d\0�gC�K�%��$���fin�lC����B�?}�� Z#�¹�;P>�e��ݚ�*�u)��%��鉏
��.j��em�qE-� X������w�@�A��WSq�:,:]:�7��V'+Em�l��1�'\0��&hE����1�3���.�+�x5�:\�����%#!"��0��:�֯z!o��<�7�MzS�͒�h�����I�3�4n_�kǹ�9�Ӻ����	�� �E�FC���`� fY��^��㷒3 ��X$�7�T�\J��ᚷ��Zd�(��zD�����c�6!ׅP��O�nL,���A�n�D�˙�S�<.��8^ԑ�ɷւ�5B@뛔];���[;���B����f��[K��E��0�oM/ψtټ���O���υB