XlxV64EB    2284     a806�a���;�m�,��o�f���?�.ļ�����p>*�C>�
 �z�P�k���ǫ�#2p�M�ϩ���`R���l.�D����˵"[.� ǩ+ҏ��`��=B-Tz��P��gUq͞IC���"^�Ky���| )������#8%eelYfcDs�aM{�26-�� ���;��vi��ku��
��f�������!4Ň��K$14�P-�7b����#wB0[[�p�1�f�CZ"���.�2���H�B���oU@��eS����wM���I����WN�K������"�%�̩����GY�\U�$�h'�9W(|���Q������a�.�Oτ澬�ߩC�ͱ��X��X:�"ָ��P��O�ZG�p���&6�a��H/m��� �Dbߒu�0[�c-�"Gԩ暩5xG��]�j��Y
1b�<�޾�k\U�*��PACR��Qkp7ٜ����ff�����N��D�[6	��4`������
�W�ӿK'��e�^�C��f��d�_�=�P�ߒi�D+_\���M����06c�OxY���DG�E!�B�%�m��Rw�����9U����KM3n���J��>�޼��f5�(�.�?�u�e�ˏ���{�Уa!(�̼u�
D�Q�@�w�ڲ*i��׻4���dO�ډ����:�̵��'�7Sp�zץ�{����xͰ�\�a-͙���3ŀΑ3���P��IF�����hs�O^�$N�p���܋�U*J�[�� ��6Ǹ��ǟ�hF��=��y���P�{�$��ݙu���J�g�Zk��fX�?���Q�#����,\��cM$�"��?S^��KF�Z)b#�>&M�]?�l7�bIl8j~Z��]Bʙ����F-nS;~�A��9�@���Y��%'Uߗ�[����ʛ0?�ʵ$���O3�� `�
)��v���r��YNOd�؟�gQp�W��a�~�E��Ol4�L��Iɰeл)�������n�����$W&Rb�贘aۤ�q�T4ޞ��W-���$X�4��go�Ͻ�'w
ى� p��G�Q[���t����6�p��P�-��џ�[��a㱸�B2��%T	��Z�$����4���=�W�xtЃ;���?����������*G�2s�r+�ϕ��C�r�'G˜�E�ZF�(���B׺�pq��I�mUI�HSK:3f��ko4��68���/֏���\���7X�p�˱(u���B$������|����׿�R�F�Ftw��t}�**!���e3���{\���(5la(�01�>9��h��ًbh�s݊Ӳ��c(+j�7����DI`�I
Dy��ŎY��	8�/��-�O�GiE�q!6�4ۏ��M��N6�f�{{z�K�����S�r�%a�,A"�G{c����%�P�+����օ�9��[~���i�L�_��0�a.OIՠZ�R�)��)b�=�_�bn[-t��|��J��#&�H��0�n�א�h����#g�D��ڠa˕g2���;@�TR���@���Jvpǹs,���3�v��x%�
`���I��:p����BP �(E�rq9n��8��[�ig�QeZ�_a1`�� [��9���mmk$-��r)��_�%9s
�3��N��r�'���V�`�t���_��@��y����T�r�&6��l*ɩ����FtBx�k�\�-xCC	U:Գ����¡���>�*� f6�@�Gc�`�	�ۅ�\'6�@'������a�v��ۦ²�{�D��WCy]�u���Q���R�Qs)4�gm�6�<�<�,ja"<Î����d�m����b3Q�wZ�`�\��R�A\��4l�y�o$Vk�)Rr���M2��@�6A�p�YU_��Մ,�E�)w����U��ս0\ C��D��ݡ�F]m�ƪ� ��הUd8��A����On�+oiV��ε��r�.�b`���t1�x����&�Ң�.�5n�O
��_jQ��c�
�W�����	O�f��Ye��ݪj�/v�l��"jh���qr�D��5}:�r$�~R����𦧲w5�H�_�~��=�D�c�Nۀ��p����&B�hKʬ��ğ�w�ޝ�*.w	uw^��=bz>��꽵k�
c���~C<,oH��c���Uի	p�KWU�8���mƋ�D\�ݺ��F�s��lg�i�{a%��;>�M���RV��x���Tmθ	b�]��ʉ�"b{&����z��0����-c3����� �N4��UO�6�h�8ݫ��EEN���+��kUe%���@��ɤ�a�oUl�U�������Lݟu��Y��-_����Y,�	<\�V��Mx�mh"��eg)��C_hm�{�Ɨ ÷�����<╏����b=g>F ���+~+R��Zz�z5*^�-w��r�,c�U�-���0"V�����@ك\�U��ׁ����#��RNϨ�x�*������D����x��EK�]�=���w��z��h��`�G��GQTi[�{�-V�QA�}h�Ҁ�AGR�4z��������>R��I�b��*����$�Y��3�̖�w-��,��^j\y��H_���5��|�>�z�)LBI� [��El�'䏊����9��j�<1�