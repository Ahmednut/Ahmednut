--------------------------------------------------------------------------------
--
--    ****                              *
--   ******                            ***
--   *******                           ****
--   ********    ****  ****     **** *********    ******* ****    ***********
--   *********   ****  ****     **** *********  **************  *************
--   **** *****  ****  ****     ****   ****    *****    ****** *****     ****
--   ****  ***** ****  ****     ****   ****   *****      ****  ****      ****
--  ****    *********  ****     ****   ****   ****       ****  ****      ****
--  ****     ********  ****    *****  ****    *****     *****  ****      ****
--  ****      ******   ***** ******   *****    ****** *******  ****** *******
--  ****        ****   ************    ******   *************   *************
--  ****         ***     ****  ****     ****      *****  ****     *****  ****
--                                                                       ****
--          I N N O V A T I O N  T O D A Y  F O R  T O M M O R O W       ****
--                                                                        ***
--
--------------------------------------------------------------------------------
-- File        : lyt_ind_ch_reg_p.vhd
--------------------------------------------------------------------------------
-- Description : Package to indirect channel register
--------------------------------------------------------------------------------
-- Copyright (c) 2014 Nutaq inc.
--------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;

package lyt_type_p is

  type array8_v32_t is array(7 downto 0) of std_logic_vector(31 downto 0);
  type array8_v64_t is array(7 downto 0) of std_logic_vector(63 downto 0);
  type array8_v16_t is array(7 downto 0) of std_logic_vector(15 downto 0);
  type array8_v9_t is array(7 downto 0) of std_logic_vector(8 downto 0);

end lyt_type_p;


package body lyt_type_p is

end lyt_type_p;