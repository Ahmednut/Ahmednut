XlxV64EB    1ad0     9e0�͒�6fxf�'n�mw�V�g��K/Z�&~iqo0Vr9L���Z~f��=�d����{�����w]�vZ����u�_Ϛk���殬>�D��|��p$F�ԥ�C&�H��j�� �Am���*��)�a������%_2�pWͿ��jEK�~r�H���,)�a�aF��@�h�?�����>��v���'A)��Il���G� �p�#����
6yP9o6B��_s���ƜY���v���E#2H��5x�N�����>�3 u��6d�
O�z�6�M�g':F�%0�f���_��`�U�h	������ޱ}��o�����˯6���S<���G�֊��}
�8��1��3ⴍ��64����8R�S�����ɴ\N�e�Xx�&U��$�Iz��3�����.�Ԩ ��u��N�Q'�Dd��L��X�u*��6��p���Yٕж:	���*�yagI���>c#�"�L��)g\\%�y*!,��XZTS�տ	-nԇe*�+|!��V7)k�����炝GŝGB�.}�9�K�������#O�<�Y�-�8�囁��:#"�;�Zx���gC��C�Q��P��}�$?�0ѴH���~`�Xs�]�<�$�"�\�8^�`yS�O�C�� FQ�y�n������@(��l��H�^�HUD8P{��ų�F:�o9h�I�FP*�#z;_Yt�9��bѩ/��7�!��9��	z�EX�Q���}�:��Ł���~w|0�ܗ�X	��l.�$�d��ayN��b}	x�ģ��y/L��{[��,%&9�A�KԍA:u֓z�5���� >f���;m-�^ ���}6b���5z�f�������{�30�C�*b�����~�g���-sqg���Y�<���`Y�Bz>"-<wi̴���8d�nkTK�z1����~���ka?P]p���Jj�A^�s���@�"�Q�Z`ǫ4	�'����q�k/�ƴ��gϳ%{V�rݱ�*M�y)&C�-�����b=�6�G�5z�/Q���:"�5�"�'�`�H�K����0#Tds�_?-�Є���x9��?W}����ϼV�^�]�P��>�L�� E�d9�ƞ/�_�ޅ����O�e6� �}�A����%���'V�C�O=\��WM!=��*D��\�);����3$hy��;�B}Q ۗ��+sD��QӠjF�{P�8��E���/�k,��ﬔeE��k��	�c���(����� ԥ�0�5�Dv��5X ��u� A����QmUҡ��G��}���U��n��"���cR�27w���wW�<^�����勑��V���ɕ5Tl��B�H͘ù�
<"T�p{�`XB��;��ER���B��,�O�#��d����Ē�۬���USy�P�L:������'is�ďE)��	P⼗Q����Nw!Gl�;�Q���jBl�$��Z�������4��ĸ|d$�o�ㅜ�ט���d:��?"X��W�6���=V���h�����Kml�1����ʀ]�J�b��w��{���xPP3O�VL�1�L�-�[�z<ٶ� �hb�̄4�5�A	�^G<߼�i��@��x�F֪��'���oF-���`�L\�f�.h\m��#��Z����LuA?׶��I�'|��-[l��}���{��.d��_Ț]�����;8h[y�[ќU�"�;���}?���Mq�~�ǜ�A�}����pn�/�(��A���G�&�^���>_iXZ���>E頯��H�yf��b�G�Vbfe´�7�s�`�wF�af�Ӝ)���z��r]+D�d��LZN�J�^�5׻3�J7$��ue$����S�����ŠL�� b<E�'A�8NO�6���~�_{6X����8�/�ܽD����b2�.��i3
a`�mp���ݓ���ґ�wM�r���ň���#ƛ��K�AJ��68R�j_ge��IW�nr���t`�"�oAy��؆�M[p��|c!�˝A�6й�~2og��HJ�;c赗�xZ������Z��=�%B�'(٧�չ�Z�<��ƫ~]�[ ��� Ym���gߎ��0cb�Y!k�f2?/L�=:�]X���	���{'����D�ԏGs=T��W3>6�!��v�3y��Q�6� nl�����&Q�0��~�ῇߌ9BMm��Z��m}g:��w�u�M��#�x8g!fe��T���Z����#o�x\���b^�J<=�f��)/ :��VA�N����Un��b�^�&��P�4<Q3}J[�x��"%���L��qVV��+��I*d�3����=�]�����'
���hF�aNK��k��V��yn�Uۍ�0)w��ُ�u��:$�R�pFɯ"��՚�$�i����-=�l�ם��ugԕ�E慊,�t.�o�5u���Pi�L��Y3�+�?�+����<��B�S؊g��$�o>ݥ�NtE
}�