XlxV64EB    1b79     9c0t�#ȉ����l�,j|��zN{e�H����\�
�`��
���c!�ۇP{�5����\�;P* $����>��QYh~�ԋ�9,��_#u�&���5�)�{�WObM�b:*���Ҿ6���JK�RY��;��$�_����Qz�<IX��?�|��eB��V����e�
��x�%�|��N}����1��CES=�[����.���n�A�Z�wxD���L�f������.���@�l�J��2
�sۯ���}��ߏ�6N�]�����b������k���C��^�f�{�Z(Q��F+�-x�C��'��{�wt*�
a=c |Yޯ�9�+�ɦ�2�O���-n�`+8Y��!�yK��k�34ɩ�o��4�w�&����� W������S�S,6}t�,��NI�\v��Y\Y�]�k:U@�1������)	S8�T"֊�'�gYuH���P����񈫉���F<D�����#Y�6��ϴ�wG �>��Qd�H���g}F2�xfo#��SX}{�d˛�����o�_m�k#�w�/NRR��p�%b�~k�����S(B�n�Rbz��M�:�[�� e��y��vM��c�[1�8m?apW���T�3A}�{����[c�V��t�M��P�z���eV"F�?p-0������m�|��MA��������]{��Xm}��'^�
��h%�c�;).�;�� �u��7����^��^�!�m�/�'��.Z����*,-S�
���� �{���e���^G8�M6j�/s���͔Głj	����jx��P���5����n�*�;1Y�R��f�0b�A#(���2�iQ����h�cԬ枴5��hH����8J�_���kX�3�j�]����t��/�١e�3�lp�����|сQ�^� �E۾|�9E3�*��w�����	� �m�u>Z?WR�8�ll�1�x\�p���I~��1,~L�,����[v���J��h���"��n@��� ��[���c��́���\?H�~5V��xפ��f���v���2�^�6UP�����s^]C.[h��9��_���?��k{Y%^]){s#���
��@�7�M6��t´^���k�:���7�Q�޲x��]pr��H�}���]@t^5V�T�B�����є���eLp���?�ƶ��?��R�`���0ߺfH��v�0޳N��5�mJiSU��ibw�R�ᢒ�/�)��u�d�8p���E��v3N�07����3�_C��M���$|��v�#Z��R���b�p�	���F�*��f\h��`p�]<|Q�0��Y�r\і��!9(3�e'&�N��Y�֯�	�&4�!��a�l*�أ'�|��ƚҦ0X�ǤĢ~�ؿ���,Yt�x�i+,4Bu�n=�����|��՛��hF�%�.#�� f�h=<G�e��)B��u�V�dg�]���y��ƅ�㴰mk�����D�ǫ�m�i���I�R�h���2�/�z�����{[�R ��X1QÏg�5٥���,mM6���]�zτ��x@����y�����n�و���6_kּ�v�+q��&'���X��\|z��g3��� N�<M@�Fn}?_k��lDR3�c�	0���\4g1��u�I5���e�
-��q �Ih�!&N}�X��G��������l
Јv�S��κ3ef�=%����,,����*'�*�kF����O�e�HĴ��|}�k�	�:h=�6�  ���!ށ�6K�`�����}���Le_��F��k;���\Q�>��̢�|�y�?5�̘��?"p�|f�bkہ�����3����6�\>s?ޒ,�k�û�� �jOuH�Ǵ�&�B��.p0��������r)�o�0�����?�;�i{/"�o ׻d=Gr��c�+^x�-�NL��k����U��H\H�w垑5�"޼Z)����[�$�fT��N`�MPPI��9���N^��a�5�x�q?އa(��:v�ry���oSZ�z3����v ���>3�"XSY���f �`�EXp:_���єr�+��㼇�jV�a���`N���̓wv"��״�Е�	���y�n"e�8����yF��P�������N��)�e)>
�C�OP*]�j �'��B�I�F-�:�V�9�� \�^�"�c��eϖ��c���Bx��)J��30�at㵴sv%m0��<2y#�b����Oј�J��ޙ���͜����1���+��q��>W=U8.����\]1NN�u ���u�a`��������������u�A����u
���)B��ᘶs춏=��f��|ƚ�,��E�i��'�W8s����B�0}]³p�{H^M��w�DKޒ77���o�t��wcI�
�B���W"�Fvr���������Í$��