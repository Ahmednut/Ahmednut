XlxV64EB    fa00    2f60�
F���^v��
1�EhtiȨ�#�חI�P|���(�*��ة����[�IZ3���l�?S.=�f-���11�'1E�d��ʸIAٞnU��<�1���0F�̱+�f4#��ˌ(ӋX�ϭ�4Ѱ�W��O�G��7y2�;bG�G�������Us�}g&��l��XD,i�=�����~��pK(jT������49&�o�g�i^ ����.��{���&;��!��w ND$�UB9)��}Հ��EdWq汞�+�t6E'PS]-�(୐���ڪ�0��� ��}Z�����5:Ϭ�ߜm��BOR稯S�UU�٤�,�����f�*��0&�o��~vߵ_v��Qv=�.^ؼ��Д�r<��(�T��.��T�e?O�� ��[�k����;��R�58��/}�����rh\>�D�5T����Z�@>���g�x4��d��}��T�6)l�R���U�c��V2&�;
^eb�^��y��"T7����f:����}�Lb4+G���V�o��j�W���J�^�ȨE�#7s�Ѳ��&�I3�s\:V56�'%�(֡CP>@�<q9�Z���+����ĵb�źUA���!Kh�E�b�8T��� s���yW<;<��hb��N6YĈf�|��ó,TJ��Km2���Ҕ8&ju �5������$ʹ�O��a�)����d�,Șp�����A���!��\ϻ������ab'�b/�����nA��;WcA���n�= ���������׷/�%u�=����k��G��tH\m^�<�L�zc����ىfE�GP%����8~�<p�o0x��D"�OyY�/w/��j����򛸄"(����h1�p���:�V6Hh���n1&�h�u�Q��a��r�1��K�oϮ��_�	y�O{��/_�cžm�����C�!k)�0��Z��z@���$$|}+��0
jQۺB`���$�r�h��]M� �h=��E��^���F'�����>pZ����i����(�^Cְv��	�����+�v�hؙ�lM5��iM/�|�]YI�Z�t�tad�d@y�,?�N��Э�ݓ�|d�~X��P�{o-5�Rk� ���|2�Y[`�������!���<�wN�ܥ��-R�6.j4�f3����G�� ċn��t�Ⱦ�Y{�t#
�����ì�4UW���eAa�(� ��Bͷ3
T��&�XH���kaVv��kXˎ}�lA��P��w�ֱ-p����j���[:��E��~��rK�aorqi�[�i{��2T#丆���˃P����1d�Nv�xV���o���x5 ��b�a�%��{��X貁��}C
�����hQ��o���چ��M�|��BVJ�����r~�;�H>n�[�Q�a��tN�����t� <ϑ����Q$k��*����L���r����\k�5�ɉ{�S΄!�s�%����I��V��[޻}���~�b�w޺�7�[�̓������~���h��x��a� �����+�QGfχx�-�aǑ��	z"0Ĭ{�#�m?�Zn����{�ɹ�Eb�ٳ��f�_՗f�C�|1{���H`��χR��� [Y�a`	��K�]%�M���aK��
�&J�J���\ەB�-�b�k�m@��RQ֭tz�i�ln�PFI���kg�y[LY��o���j�H�gU���҄?'H��{�=��6J� X>�i�7��һt4"mFJgرe�@
����k�J]��m�z]0�'&��Q�������J�fppA_o#�%�����alN�*F����i�)�d�!/ �F�����qRR�mݚ�fs�# Hԁ��;�"ٕc�r:���Q%W�8����Z8c���?�����K0y���O���V|E�c�RO�7���l��b'�1�Ό��0�8U�ء'I��i����#z����[����T�
*�|��[IS���f�[��*�����Ma��'Z"��&Cj���gQ��cphu)q!�����=����r�X�	�)���pn���
�i ���b�H6q]��r[	��͑��0��n#	Rّ�����v^�^9�DE��~9X���^Z�e�_}��$m)=Ю���WY��o �o�m������6�����}$����tic�N~5�
qæ.�ͩ�����#�<G�&���C{2Cj�/�0r����J�������pmg$,����(ŴQ[��UՆ�y#��H02̅�������K�-_G���eQ\<]��
q,(qj��d5���`�g��9,��6�������b�2��oN�'
5�\��?݋/�7(;�UB�����FB�Q�(�L���C��KShF>�p�/�cG��|�Qx|��f-VhX8_�g�'<X���F@͕����N
��ɾ�T�uC�\�6�خ���M�>����!玅ʴT�lV
5���w�(�B�i?�k1�z�D��";��́@��#��˥��f��(��	�`u�_��v ����'_e4���p����2���Xt��+]�+�)w6P�J�	��ώ�(��^�`���K�M�m�V��ƞ�˵�Z�!Ɲ*7�1iS�hA��5F�m'�aR�VN�A~��L�C�V�Wio���uF�u,�Q29Q���R��85�>�yk$�]�(IS敍f�r�W�y�	XT&��:y�s�ɺ����;��rͣ
c�֖�f���&����ܺ�����A�x>���}��A�ő��(JW���\��u�W'QHP����`;Pu�W3��:�v5�Fo��g����iQ����3��Y�)���$"N�B��{ �g�T��>	�{,#U��/���:��X:a��QW�?}͍�k��s�q�}$#��8B�oX����x�>�m��<�%X����e؏�U���s�/@Oӧ�Lp��G���ۑ��|Q3 ��
�AԼ��ޘ
d1��&��\x��zE��L�ßta�������]<�?M�<[ǔuf�?ȲI�D(@���?>_5��:8�%�0}�EĀx�S�e�c�^M�i/����P;
&�a�5���ņ#���I;����c�A�$�}+;���� r�&�ǔ�v/��g�p��!�5 �E��4B�,ǈ�$8$>čx�n�`Aį�c�3�1%��c�.�rAۙท��?X��Բ�K�p"�v_VD7�$ʠu���u$��d��\�c�9,Qxh������k��l7����w^3��&A~������g�C� 15��q���}�f(ʖ�5��<�__��ʡ��𛜉���~`U#���e�:-����Z�-a���.\�^n����N�M�.J�e"����͔k������%��#�P�g0��v#��Uߠ��6�+]Ȇ�#Q��J\�Ga������W�[��l���w������p��u��T��v�#��e@o�w�xrE��.��+��i#��.��z���>%{FnX����3)V|D�s��^x�0(�~��&����UI�yA �-?E���IԡD�o�H�Vm���2�1�27)_��~����JI�{�d���B���G_��,m�^���N��Tr�cm��̥0�
jA&�Rژ?(�~�x�Fqm+��ڒ-,��ĚKy�����j�[���Վ�N�o�%Z�_�O5��H����b�����+����eV&�*��~N�>�R��m��]��E��>Û�
\���F��Zؖ��_P���{���k�CF��NX��{:2?��/T�X�Q�;>G~�q��WVU<VF�~#���v̍Kl1}�~� Nr��r��o�1���i��[UuZ��i��*��+V\���oB�J+�����E��A<�`@XZ�8�^<���f e0��r*�0�Zߵ�K[ʤ\�5~���Ap��HVY�xY���m6,�H�x�a�p�$-d�"#|���TuM�d1/SY�セ�	J�����|aȊJ�L���4�>(/Q�9�j<��G�|�����ӵ��1.+�
�
[�;�9 2ϻJ/�yE�Z�чAg��g�ż=�dTH�W���=���r�Q����Th�&���$�p4�m�_��F.�0��>�����
7-�j,CR�U����$��4����SNf���u�\w 
2/?锆�:5kf�f�׏,?}� Y7g��gn�E�Xm�T!���t8��1'��0B�Z���Y/p�~r�͛���U��L�L^��� �
��6������S{F�it!��z��U����g'�Qn2���JS�jڌH��ܖ�����q߮���Dm��el��p�r����.>FS��:�ޠ�Lu�nF�B��X�K�&�B"����b;����y�:.�9t�͕�T���q�A��U�ޏ!�����͢=�Խ��`�T���{��C�������5K/�DJ8b{�mQ��ۭ��Ak��ˑ��\��p�n#�S�v�'��MB��YJq�9Y]�|<��X謅=��	��,]�3�65��{����ܞ�1���Зm�)ǿ:0�~��(�4pZ����|q�C����J�3��f �'��-��	��qHH�a��K���ᒥ [�����:�b�{{�D�]pz#�_�-t��zT��_4V�WF��rO�4E�%�le�Ru9�{Ȉz����b�1�<v\�'F'�ĕ\���q��ԕ٢���G"[_�~$-5\����s �7Os��@��6��$N2�ClkC�}��L,�W�1��lOi�C��dS�膒��B>�rN���ە�i��+�F�:�^�%� a�5��'��3=x��8��*�G�H�s�~��8��|��� c���9��S����0;'IT	ߐ���Ԗ��������A���2��cH����Ǖ����v����i�0n� ��{�bO����$�qS��h?�
�C����c�5��Xʴ��+��q�l�v0$��;�F������9�ʊ��[ɌҲ:A�f�ڷ���όc:2�r�r/u�� ���,�W�O�)e����e �Q6�yk���o�7/~����Lsi�UCkK��\|����5 �D �AH*Lj�윱ko�`��9W����H�ꎠI�6O��7�yJk�]4f��� �Q��]�"4 .���6 ��������� �1*����)��ZBa&�38'�I��d[�<��Et�E���أ�ε``��'[BF�Jg��|= �'�RKc �Ƃx��"b���X�,�\����{%��n�<8fH! f�"��QB�8�6��+�;L	��6���ǐck/R��B"|p"xtL��-|.�<[�t&�%sm�d;�������,`�3n�2�\�NM�݄���M#���R�PC�Bv]�ձ0k�n�as׽�%�5r7�����6kˠ�[���v4�<Fj܌gg�^܃ӗ�"F�ۂ��T�p���
�u �A�FY��ୡ7f�~6cG�I&���9��`�h��r?J��3�z�4�U3�GB.�S��s�"ER���PBl<4o�Og/�F�In9Ƴ��e�ObaO���/�����0$[�__�ԋ.���Z �[p��m�����cӈ�q��u�Na�cS�U�� >��§���kjW˧h���`\�	��-��B�J8S#���㾖~7�ص�G�>�� n���*��*J[�ak�s�_\�'���n�\,�<�,v���!�U6@��0lI��&E�|��B�)�c�]����9�uћ�^W�ʋ{�����N}������=#n�n�c6��}>�B�Es���eV{h.$P�f��N���xj�tU��Ɍ��R�Ѱ���hC�R��F�uG}g�tR��SN���px��WHT2�		� (��DW���ޏ7�r.nd��m�����r4�^zu<��R� �:@�D
�F�A��&��Xj�
\�u��3�Ҏ��y�9_��#�Ę��;��e$���٧�;�Y���t���`E��2�~j����I ��1!n!G�;�B�����o����]��C�o�Y�/���/F�j4��0���S�Ղ?L��l�WN�/��r�z\�%'�$Iސ�ϥ��X��b�5�#N�7
3����&�m�������n����Ō��Pu$,���E7ʻ��2�8���n�-�K[�ӂ�����z4G��3�>p��~����d�~��F�(�Ga���'feAS�@����Q�](c���ӹ�N'{'HT74D��,s����HKK�MGHw�if��,/WR�^_6Y>>'�v'^�M}3���ʚ&c
��z��,����X�_,%5��x���5\�5{|ع��U�z�߮��Fv��@0�y.f���Q�L��F��s��;RC�`4�1ewיA���n�� �~�$M��)dO��v-���Y�$0�,э0k�Y�������f寎���A�׫	����2�����I�q�"i:{ �K�.�u���~�Pk�o�5��B�����΄U�^hv{	LJ���a�ۏ�er��.��)��I�Yd_iN�2�S� `�A
�~�.��@ga1nc�5u,������g.^T���VӒS�C�2�f-���:�&�nV��{��Y��Xe��9�;'�I�	�G�m�o:��\��Zw�J�7����C�'�������va#V}������V���4[bo�s�NGXK��$�%̱xjI��1`%����5<(	��T��8���i�if$��Y�WLq)��j	&�[�����e�$3�u\�-�Pw-�������X�E�bMi�B+�t�ml�
������TD���p�Xx]]�ܛ�������uNt�N�3�� �#�W��*�&���r*�A;1,!s����N��^����3�딄mϜaD��+j,f"�^��.����L`�5ag���L�������>�6�I�g|����4�2"�U2iZlV�|�R��w��E;��8	����Nh�s�O���J��>��96�����AD\��#�G'���2�<��vHs���ȉ`-�'0\�Q��/��8��`�Z�T+M�<��,�^� ��V�^�o<��� ���%I��A(>�!;��$������+Ygom��תu��,j^�����3)�4���7��F�\0�	U��a_jE]���"=y.�gUS��$�d���F���)-n�<%@fW�r�ݨ���L�׊�N��Rne�������t�ƪ������E�P�w����[����O���l=�X�t�sh���^Vy~�B�T��[���/R�-�?r�<ɐ��À6�����鋈'8<�87���#'��jg��T �S`��z^�^����9�3ډOKm���.I����Z�a4�C�C�A���s�;��0��~�S|�'�O�<��ޮ�"I�_���؄��)��o�� ����G�Е�_9����#�\�~GhU$.�s��ƻ�#����p���P~�W��8F��²=r'�g��a��z��k��W6�t��#O�0����)3��*EB=y��ŉ�md�,�����Hhc��b���s�Y�)᷇�p�{��GK)Wq��'��|<�|�bBuk���N�'�`ZY�}�����7_���Ž`>��i�j�2�I�#K���!h3WC����X��yp@f�M]���7g2Mn��qg`:�yJλJ���~Ν����&H��I�����N�Jy�4���j>�����Ջ�!��u��7�v�W�-�M$�0���J�I	i�_����5��k��G=�`�O�s�j�������� o�������{Et0�53㜶ʵ��#dJ[J�:��3�,1r�f,��$��wP���VH�944+w
���<�{Ż�'��g�	'K.�7��Vtq$�i�髍�"�U��eX��	Z�;�'�
��?�/�${�b����i@n������S�ݒP3�m�Zɞ6���G5|���E��_u(��O�@	LD-ꋫ\�2�rw��	6$�����7<�'5�i�޿�p�t�P���'�<^]�`��3>����]�K���G��G靼DМZ��b�3�U�^�X<��a����l������3�ȷy����[��8�\G[�C;t�b����(������H�7)0=��ʷ�inE� d�.H��D��uWUZW{~��Ɔ6�Dr^�u�8]A�����0�r"/2��n�M��!���AN�Y �z64T;�5P/�d،~I�hykI �fOS$%l�C�,閚"C�|�|m�,I`�_}�I��(B�����Y����&3�ݚ�n���2���*��Q+���3`�V���p�L�vjݫ��8SHRn0sb����u��HW�����6����R��CS�<�,lA��'߳�&;&H_I�D_�yX��0&��������i�ׂE�8E�P27G���\�J��I-)k2�c�W,���?CJW������d]�50wT�d�5��IÇ�t�h���|"��JK/A� �Y�a��z��Cs�oN�H$�@��6jG4ř��n��v�W�C\��r��t
�pT!łu�c;o�(��2�̀4���i�!����a�P�����{\aƫ!b��r��i�e%�� V�1���8�� ��R�Aٞ�KZr�����Lfp]�9�c!įW��]h�����R�^=�p(�-�~����ý�%�����͒��D.��"[N�uP|�G��1]���ɋ���#D{��AQa`��z� V ��(�q�pz��,\ {��|H�ٖN�KG��2�T�ܨ��},;>� g��N�����g���|�ёC����i�����܁�@��M"��lJ�PQI���[��V���� S3�H�9�C&��.UO>��6âG����1��Z�X�B^N���8Og7G��A�%C�޳�uR�����\hm��dt�
-�Y�n�#�X���3E��2th �Ne���."���m�wk�5 ��T�g�Ȭ�C�$����"���x��N:@:�����oȝ�2��]ρz3�?�*��M�ǔ>_��~]J[�l�\�fu�`���crL�y�H��9`NN����"���={m�D�~��lCh���hY��2��E��"��7�l`�Uy�H`�HU7�ƴv �Aw��J�*[BM��#CN�w�g���2Z�Αf��O���_���)$uY�7s5 j遏c\�w-MOG��3E�5v�Q]مU:M�0)='99�o�����HlKGyhA[b��F�y���	�Gl.Q��`�\��7giL,��l��AO3T�c��'��$��mq#V-�i��ȕ��\��g���(Opcݕ���wkYU��J�M�>ÌbV���w`���X����zVe����en��𳸿s�G�2����j��gwr�KN�׎2ǋ`��E�'����;Ɵ��p0i�á��%*�hj�W>+��Q��ő��0L����j���{�x���'b߷����v��:W$,�k��w6X%DK�4S8�(�\�W�+v�Ĺou�y����1N��*?��gc��a��6���
K��>pmo#��B�D���pL�	l�y��w��ѧ6~��*˅Q{����T`��-m�?G��y&�B@d�@��HƟm:�i���&�K�Y%�^	*�fw;��2,��-25&�A
kՆ�v9صbW��f{*]m\n4&�qz��_�m�s�8*�<Y��FNUN��"B�S�Ϙ�B�KZ갌�?]���3 u��J��:�V�1�)��]�R��;]�p��;�>3�U��f/H�c=���N#h�1)�����.;�/��qjZԫ^�c"���������p2c�xmb��zJ��:4@��w@�������(��u=�1��7)'�骣Ĩ.΋�1�)#\j�l�mÀ[���W�M��c�~�ݷ�E,V{���nء�\�qB�uQ-�7gC-�-�Φ�yZ2(�}:������h��s:�,�ܣgn��bz{p�'S Vj�Ԅ=��hC��O�>���nR��W�򖯒� �'�!��D�C&	IE��0n�_P&���Ϋ>*��I*�"�`�gv#��zŃE�l�8��4c( ՙĄf��*�m��"j�t�K�iy�p)b�����_�o�ϟbkU�\+���2��Ⱥ~�{Zc�����<��7hIM�A�-ͪ��c�#0��h?���������c�8\�ߜ�O�HT�\�.c��s��j$ں�i��6��gr���=<�T2ZĲMU�D.*�@���NΝD'�t�=�k��pm�԰B�d� <�6�]�
,2J*QI�}Ku���3IQ�xa�rgn/e3_�ҩV8�= J�T��%���m�	�=�s��}���&�+PKR@ê�I�"��1q���9f�a@��&y��	�I~@�x�,��v+��w��X	�9̿R�z�������X~`�I��ٟң�Y��O����T��z�5�*^���Ea+2�pt��m^8��a�i�����M�m�O��_^��ݼd�sTq-�'��b�J�Y�$ w\�[�U�}�"�_�񜛚l�V�q�D|`^�7ĩ�1�F��8��?k�8��"�s�
���l�Z�*��W��� e4��{�&��{�V$d��`�N�֊0�i =�������5�V:��*�Kک�@1O�ۍ�#(�K�C�����T�3�i+�r�ʼ��ň&UN���c@f�bi��%���1���b�cJ6�����9�5�x'Gy��I����>8�bk���Ѐ<u)�tisi
����!��Rn�q��c�6)�����f0B�
��)�U&yt�W�c(RD;��.(^$�V$|�y�4E�d�B�P����jڠ유��d��"�l �(��b�������8���$Õ��&mf`�b�w�U��إ�"+\�G�P�U�Cb��=���F�Q����d�����wXK�r����qB�wq�9�K�^c�s�g�Ϟ���FhO,�VMJj	#��	L��b����X��φ<\�	���.3t,gƟ��^���}Hy�4�� �!�P�V"���u��
^VW��V!���㧟�FQ��@�{M�Þ��%͋�U�@Um�s�VL���QT�D��Q�!���zp]�~*�9�
�v�DR���5����>"�+iL�#7^�s�Q�)!��I��;k��7��~�i\e�6��� F�V|<Z��-����
*C�Q	�6�f����݆3���'�����mo�(�V������C׬���n��bm'�N�p}s5������q�M�Ƨ9�'�ډ������B�}Y�D� ����v�@�Z��;L��b���*�1�eNQ
��y��]��_�)\v*��:���&mrj�Ʀ��L��+���#?Gw�f����ًO#tܻV$���%���#j�V�����.���6P(|� ��l��v�#��r���E2�(9w(5��H�q�G�!��
RH3E�{��o?���SD���͏����F�i"���>I�L�=�ݥ%�	��9�F	˯�7��)'����#�-Zp�%�&�[�e�����@����ժ|/%��-o��S��=[�+����Ł}MĀ�&H�~'`NXhc�߯E��\��kQ��;g(�'�b��/fCn�N��]d��� X�A妚=�$�h���0����S�t��Ψ�7�Փ9��r�x)tvj�c�<����-�;�}��a���Y��fU����Ō9�,�H�I���Q��L�*{3�8��g^����\�4_{�:�Nx��d�ɬ�H�-���:i�J�フ�twPT��S����>��Q�Ӎ���֯gsʥ>������֐՞4^��u/w�^/��.e�G:��2\52��P���O��F ,��o9p��gW�騖�����҉^���?�O!_�І?�/��cZar�z��|	��:E����'���zFʛʕ.��&���#RyXlxV64EB    7b70    1910�7�`gwEXe�\������X��E������>y�0!�>u�unB�Ǟn���?.x��)eYB4�h�3��r��2��p����CΟL���)O�H�x8���s��X�KE��wԿpq=6�E��tY~�->ؓ�E��7��*j��W>�u;�ڡ�B.�B�ʥrW�!���a�W"wO��^.�Nk!����MMNl�&��n�����6�k���^1� h^������w��=�Zrz�E�M���ˤl�'�r�F�`_3��,S���W<���N�Ք��55J$!�a�$,Zhi�gN`�V�ڞ]�B���"��1����f��2ZM��]Q�[F����L���Mfd�W������%��ͣ.���.Ek��Дĩw�A�(Qv��u����/��&���<Do�AP}򬩿��CB�X�^|��jGtYW?i]�2��B��c���ʀ��D�d�Mt�}�Ә�l7��3Y�<r)�Y��3Y�i1��2���!�dT.����@b��Pp�d�� s���+XXX����#k�A�����YO��t`O!k��0T
�ܩ�y�WD܍���ۻ��d�M��em�O�v��Ի��͒m�M�u�GE6��Mg�O���j�A_���~���	���j���\�}[�����s���Pa�&������O��~v��Ps9-��5����j��ea�"��;��׎8����;Zu��P�q|,��B^�Z��] _J�(�\2�:��.g���Zi��1����)d�e$�g�v9���[)㽟pk�	�E��.v��CN�ɱ@������Å��<�j5I�i�BT8Vb?��(��kD'�g���`K��I�p�4����?c����JU�!�,���#�k�M���8��o^��|�]� ��	�\��n�Wr��j�
չ��_����G�'?�%t�eϺ����/�sU�`bx��p����iɖ2w!ǥ����K�B���CIi�1.���*d���H�߁��h�ꛆ�/$�k=��.n1���
-Z7>��p ��urϮ&/Y�b�1t��r�����ʾ�Y)nsvqhQ����2��/S&���^\� ��c�~��J�����km�Er�(|��gS�C���������w��k��'r`Y�K�:'ĞKÆ.4i� o��MhD���(aCd��)b��j������F��rjڳ��I�6�˫��ÊX�2��g��̀_�:�� B���꿹�mwЪD�'e���ӕ�A mG���p�J�;�/����O��7�H�b��`���������F�Zq
"8����)#a�o�_Ǩ��f��%B�c�J�;�ʊe���vջ��`6�%��W��̢�7M����o��5q~`E�ӓ��"Bw�Pҕ4:X@����UO��W��r��ٵ�Uo��>��k����Iŋ��������]T���YRh�)�$���F��K�\w�y�{����Y�F�� �LF}�33N��N���]��=�6v�1w@%�����0~Ȣ-��Kʠ�(JX�����.J*�Q%�j�XY�B�V:�&���zر���MjcP>,�A�(�rOAB���֒Z��s��*ۗ��3�(��$�x����Qx�O����윊K�I�f#�c�46�/�m�HP{�����X�@e�z�}R����]�l�ǻ�;y�:@��nQ���q�x��k��F�r�e)�b�	�'Q�Pf�-O�_J)��+/zC�D�K�zR�����:��r��\�j�*|�M��K�Gw*��h�@��%jEi��Y1U૓�y)�J�@nk���:rA9�	�y��ƪN�WX]�W���r#��QYXu�B�(0Ƙ�(�� H��2�6k6͵`NZ�,"�t��S8�?K�9��~7>��vp��;��A�R��C�w�1}	��Pn�4b�j�A�x�d��1�1/^���Q�F�?^����tR�dd�P*c��2(`�
$@�U����h����{.s����n��g��:9u��A�`�-��^a@2� ��h��&��v��k�T�!���짳gc��r}���������ը�h_h+(����?~D[X����ԃ�+�E�-S�Py�6�L�t3,*8��q�P��Y��phf{�fSg��gxb�W��n�4�8ՌUZ�Z�i#��?e5F��X}fV����r���v2�nŻj�G��݀ �1�m�O�����Q;�h������J�\���u^�j-����QΖXV+�'SsV����W�Y�r>Ʌo}�'_���`��`��X��@׬%���*��nE�"�;������;��K�e��G$iAo�MҴ�,���KI,,	n��@t�]D�O�}���Y�E���8�.�P�*���ß�o}��(�|�DdR�� w�č�Y\$)�;�Qr&�1�	�cvߒ>�z��}\ �R[���YX�5�e0i˶��|}��[�Ue�]��G����D�DS�I&��{0(��M��͘ %��zk����R�^Ų�TWOO/E'�t�\�l��J��ק\#`[���N��(Rp}Oޞ4�V@��vc���~�t���P�'�\
�!��F�����d!v�uyE����|��K$�@Mo�`��*�>g,��m��=�=�-�����F�e��v���M��	o���F	4c�'�n�0��ډ�q��V$�N^׼��V�V�8�z���U��p`]$-4�L�+Е�"�2��_�=��5��N�G�@�����~�K0���@�۪!k7��>���.���`I44���.��" Nl�By��� �	/:�*^��%"Z�x@�qq
�h"�[�R�aV���tb8;�ݨ��=	g����8͌:v�pUq�S��3��XhJ��R�H?>�0�8���  Z�)���'�Ɍ�3'�zsN/s�Nr���>鳞��E�_���e�@�3�;
�~�E5�U��P)<I��E�[�v�YE�q>�Sl��A�,�^4�d]�Xs��Y;Q��ER��;�e�U��!���~�K�.�Q!�V���9�1T��M ��o��lor��""�k	�p���X�}�>o���U��S���N�4����e<�K~'Ѥ;x���S垭"M��T�{�'���E
'�0��48�XS���9�����#K4�Q<�f�8�fG���P��.��zy>AlN�F����4!���d�e݆/���C�Z#��x�b��@Wr{R�1���	��S�nhA����� ak����N���f=*t~��"@�j�n�����==%ʞ��|�t�n���S�$��um�dlv/O��	��)�x��X�� �Ti��B�uc��X]^�9yUt�v�)w�+Ir�D9����m5�cw�q�x �s�8�_��[L:�a�[NB���R�T�3
|_i���3�J���c1�O������kcB��L�6rL͘q1�{OG�B�|3����JP�Z���:_��4�I��nݟ`����,Y<:'���i���<7ّ8�!�LF��o	�b��'������ �|B��"��O�ˢ���H}��ڋ���Ÿ%����J�X*����#@6��T����Ґ%�:Y��&���&[�o���=o\�W�T�\�h���w����v�-���ؤj����e�O[�e��l�XgA�C���2�ї���_6���8�ހw�4}��Į�HBe�g�ǫ{�wlv�o����4m��+�l*Zҽ���z큸�H�^�ڈ��G����I�S�AX�[��YQ�7�▭�F��!_!�������2��U2��;�}ߚ*tIom�>�9� ��ՏFJ=#���#��N�]��ΰ�zt�_N*�w��7��"����jr�� �"��Xq]z�6�<����2iu"K�ѥJD k��GR|���M�i���"�N#"t�9��T�(ަ��t+Q�+�j���N��J��s�>��)��Lu�}�z���3g~�6Q�U2�'O�G���?k<�=T?������>u��ݺ���<-XUޖ����u�J�&��1�C�T�Q�i�G���K�l�uf#N�ؒGW+�� [(��ok�R:�5 hݰw��g�F���|��:I�9:�!�!�@:p�4-,�WQ�Ba_�BZA��f���׿�IXH��sX_Z'�nے��an	D��-�pꡌ��x5]�]����[`;��� 9l+^���v�g��ݢZ%������H�u@"3��Mځ����!F��9�"�#���a#	cQʅ%R�'�&�	ul5X!ׄ��urA~kL��BfI��t�:���mTE��4KpE�S�)~�
J�fy�"�O�@\��z� �=�?�_ �Dt/l���c��I�����H����J�KDm����+d�K� �pƍ2���=cH����O� y��?H
C����F&��h��㱃��N��J�KԺ.q,�뺷p��㗫�_Ī�kXb݂�������3,���'/�4��T5r[>l�ȁOYc{L^k"5KQ��I��pZ��4�%Ѓ[����' :��A4������,�,<��aw���a��d'�ގG��[��%��Fm�+v�&$XOx��g��ǣ]��Ӟ���w����;��g�"c�*iu�w�H/s�HO'g�r�����Ƀ���@���E��R}�k��gK�',E��.c�V���զ�u.�eL,`IT�^��T��'*7�`��M	���̋z�ݬ�!��`����ؐ,ȃ���lܭ���,G�`6�Ew�^����2�d�ųYR��MQ�߷���� �n�� �.��Dr#��o����&�X|fg��dN�-N^�U�#�S\F��﫲�����*QR���(��(�a�4��+n�{Q�#����(�eۮ;F����i�dP�@\˿��*�M��9e1m�79K
iY�T뼑�73�#�����Y$mh���bG�{L%��sA7C���)͝oOw3�V9�j ��;���J��������`�������EbɇSڬko�(���>�,3�}�!�ayX���"Tՙ|��@���AM����q�=Y���{�΃F�^Vc?Av�s�d<�\&H���Ԁ�+�ݡ��vf*0PeO�������P�M�R"��{��-&���|1�3�"Y�d�­�ӊ���q٪�񋁋oc|Iy�3y�A��o�6Jj�o�p��^8e��Y��$�"��R̨���M�\[/Peͷ�����c9s��K0�	y5���>��r@�������L,|4S9�~,Ґ]V��xj���2_�5Ftb*#֪��1[�8�A#��ba����?��ϫg�����f>f��V0�H�QU7C��?���ͬ��j�K�si"w�e���/�&��m�� )�nh4 �����l�][<��δ����N�d�t���@"��Ej9k+.~l�'��+9�������]������Z2��2J�1�����a&�(�9�� ���[K=���Uu�k�>����?C����h��?8�[��Q�Ć)1�MŻȊ�T���s����h�o�򝭧Q�P�&�K��d�ѵJ��.o5M����"k����2 �0eq��oc�����қx՟�.675��1Y3u�t��R��r`;"u���'����%K��h8��k�ǪS�50o;L�W�m�{>�u�nA���VkQv��՗��5m�_�=�-
��'��v����?(��|H�/��>r������WD7�<T��K���}�;������y��֔���|�٥1qW��7[8���2���o���\8�K)p���fA\OC�%��d�q����F��x��"�ј���H7Գc��~;�rdj{b��9Hfl�PQ>ˍ[P@|O��UV����Wהu�a�s�\�$���ժ�R�����Z_���-ԙ�~Sa��`���)#ŋ����Z܋��w*�ҡ�Gy�t����ɛ�o�2ǜX����H"���y՟R�Z��z:q�m)L+:�Ӊ�`�_��!$���K,0��R��̲����)X�����ENx��h��$^iu	ޤ�(R�~���)$=����fa
�����?�[�A�ys������X�3����g��	u�UE^�L��O�&Qϔ��H�@�|ʱrk���^�~m�G������&�#����Y�ٗJ���_D������?������{���_�SF��7��4�t��C��Uy�P�o���Ăʰ �����F�N����ۉ)��ia����D3Q����Ή�X����+�U�HZBkI�?_