XlxV64EB    31f9     dd0X	/���Hl0h=d<��-���߱$V�j{��]췰!T�˜��|����7�9����d�,���O�ؓ�?o9�d�iwI�����D�Cܡ�Zs���:�D��wbC�������\����-H����rx��AR�������h�	�!(8�Reo�e)}��J��)~q�uU��<fp����D���֒����"�ζX sk}�m|;1����j^�5�r� x�_"!ŷnS\g��P�B$�QT�	x��w0w��`�&�Ps!M�f��ٳ]�F��k�<Vᨔݠɓ���nac�GX�|�ԝ�9ܶ�H�֣�K�{C,���^�G+�������+p`[�(�1G����E����2���N��!\P��^FNg���E�W�DOǀP�B����7��V`T0Ӧ.��e��@Σ�����?�Jdt�3����Z�MƱǉ�Bf�B�^*�ӡ�w� � ��H�]ʇ瘚�M��/�}r�t��p(����e�l(�3�w�>����uX�Q�\zޥk�5t�T�{X�̨d���cl��m���Vi�'�W?�s�.��:�<Qe��Eo˂����䢎~��f9.�aI����l�̎T��t⥣<DeG�.3��κ�cB��\�|P������$������	נ���";��H.0���Ni�:׉��*i�o��8���x� �l_v:]!�D�\Ӭ#"3�1�"Q���O\	���]��ô���#�O�f��ɘ����5�t �۩I�i�w/�u�!����U��:�G�W,�@i���me��F振 yG������v�k�>4�M�f90I�,?QW�:6�V}6�W^� _EE�^h�F�=օ v\�Y�r�kK�~�~J�ح�� X��<Q4  m�z���&�����zo���q��S���z"�X*�w������Y��/f��\��H�X2�HH��7]�닽���a?l��I$4�rt@6��Ū��"�_���(q5� ��T��_�1����o:�*r2,���YC�}s�~��s����J��&Mڃ�ɛA�B��̜���q\-�y�T9��cUj����S�l���ᓐu��D]�~5mA� ����/�f=�E<�È�8++���k��1vn;�<*��~�.�[6_#��ƫ}t�¼�V�Y���N�����4Ӫ]M������#��ߛ,�tgsj����%� $��z�����	������uz�:�cu@���7l5��K����Z��x���kt�Đg��>L��7�,�[z��x~<-��?6���#�)fOF�]��ݕiB����c�ݲu��`�O`
e���ٛ[�6O�`��M
���1C��7f'�:W�wp#��IA�Y����,�B�c5ݥ�=f��d:����/�1��2�PXT<���0�֊@���earUM|(��0N�:ģD��{�ب��
9�FO�?�^�^��B�2KG�q*��a�o+��gŏz�'��l�k_��x��5�ԣ��}����0:��[	�X�_a�he����i?S��q� ���x��*EQR봵ŏI��Ց�2����aC8mQ�E9��4�0b�]����Ӣ�Up|�7^��x��?�Hko��� r�����lY[؋�r4��L��C��wi���쮳����=���<9� XXs���V�ʰ_(Ԧ&�0ʗ�%��>�@)�����i�g��h%�UJ�� 3Ϸ��T�#ԆP����n���l�g��c���L�m�~v�L�^c��>�nOտ#��vƇ.���j���`F��(O��`Wn-�~�ب<�9NP/"���f�~k���hQ�і)�n��Fo��y��)�/�2���Lo&A-��D.a1��VP���䖋�L�T)���T����ňZ�k�5�����%лI��3po&!�r��6���V�Ӣ�Ewa*���T���f���P�F_P���/ƖjZk�V`EU�y�y�٠JƄ��v#8f-ZT�=��Բ�u\v"�t/��L
���5ٟ��^���n�j�,� q�p���h���Nar��"�A&d�+�vl��u:��%)=6�-�P)�K'��HX�gs�,�u�z���4���w<�-e�o����%<]�.o�ϟ���:�\MM���ʪ�����X�<�xS >�pݗ�@!b��f��+~�E���ts:��c �
m�m9s���7�q���WFM~+����B!|���I�o��1�4�fׄ����ēαIO6����"��cj�Q�9��p[���	>m��B� %r>y���ÇҴ��(X�|���5eA�jm����>�s̶�.Iٞ..w;k0��Sbљ�(�� VX4��+�?��j�4���CO+Z��4�ʝ�k�]#c�^���A
Z2��(�p�ư��%ޔTxQ��TJcS!��VȺ�ȶ����Kx|6��Y�4\B���ɝQ�Z\�<��y�:$�O��cD��Vj(׭���9(*:�;W���r�k���MFv�C1�2+�:α{�GY ��m!����
{�o����ƭJ��u��w�(6�5,�: �V��e�,�\��@+��VM[[�Aǉ�Z|V N�k�6� � !:I\��I�l��,��%�W7������ߓ���=�M�X+��;����ŋ��c�aKI�Pp��s����X���P���*�_4�����ByJƝL O���s;)^Cm�t$�>Ҳ�&�y
�W�U�P��`�����OU͍$¬	QÊ��uA�?
���*sw 0�R��;u�a�;b�w�p.c4�F�D�VF�50�ۤ����mr�5e̟5�]�`v̅����*�u�C-�7QH	�	�̏Jۈ��	N�����i=��pCF6}x�ӜG��G�+	>�-��ϛ��sy��?�X�n�	PrB&�F\�:�����(;^�y��h���G�Y}X���E*���k�F�:�<��9Z-�qܶCsd��l�,�?K����/�`J%��q�'��|��(%,f����tOB�^�@�|;y*��@��ށw������M�{�Ȫ�~Ȓ�c�ʡ���CN�W޽/D[b��}) P�uHN4�ϵ�&@�����;��K5�$�|�qNJ����+U>����I�Ӷ�pE�V�(@�<;���hO��L1E���d�~n���I9�C+?E�M���Y�t`�I��
���E�-�~V��>ŭ�)�o��=8%t�W�^�k������(��kc�؇G����
�Z��m��BCQ ���kv�Nk�����	�\�/���ǎ����P��[$�J�G�Y���U �|�8���7�Bфhہ��h�r�e`x�hdASA'���S�'��ĸ�X�d����I��+�"�ۖ����;t߳2҅9�K�X:�0���j��޸������$95D:|�Q�t����1��|���a���w�u�%��$��q��1ħ�9���`�NC��{3o�����