XlxV64EB    970b    1dc0�D�k��w�Ro{Ş��v]QM���	�g:�Գ��~,�6\�@�VGP^&ŰUiU�3���?�^r~^���~4g���U�K�3H�K�� �T[����\aY5�jͿ��q���_�	�I�mI����}���xk�V2(&^�ew�(�A��Y���#�N˗ˤ�Ë;n�b�bQ,T��$n�zWP!`{}e�^JYe8��S���f��=�܌��'`�?�5��{�=a\��W�OSH9��Q���y�Oݩ^(��!�8�Q�n滳
ٔ�KC���Z^�|+�$)�Z`^	d1U;�*B������'V�I���zؘr�j�� R��.a�2ww�I
v��R�ݍu��>���a�al���Og��1=RsH�	��#�:~EOH���⭕O�ء{����I�]����d�T���Y��$	Ͳ����ޗm��i�'���`�p��/��THѝ�U�ǫ/q&�O��s��&�D�/]�R�遑�y�ZN����0+��Ί&����<K��F�K7����֩��DX~m��^z�b[Y�GۥR�h8�/�GŪB�[k'6�`eb,�[�1��,���"��r���v�+��h����7�d��W���Lƺ������9m�.Z[1F(|�<EP+���ă[�|d�u�ÒQ�s>��PlhB�[���]�k���hU\>�?Ѝ���\v����O饧wI)��8��X	��<�9����$��f6����e^�bm��H�J���F�p��*E6%���w��8]�ߒ9
��������4k�B��րm��f��,P�;�N�p�H�`���/Mz�2��?��׷d
����)?Q8 V@ic��V#�ͮP���PK�i&�o�k ����a�@#��y��ÖU`���#���zCc��`	J!�Az��#%�K��fO�;�8��h�2L�;7�t��N卵s�X�O&�ۚ_`EIO)Ni�v�έ�9�Q���ɲy��vc�8��i�vǕE�(���m��b��]*'Ր?qx�}�?�$����˿{כ#�X%d�{�T�H���,�,�J|�~8d=��
�TX����A��t��k��j�|Uf[_AX��e������ߖUM�^LlZS����-�aH�T��A5�(FQ��{��]���/���s\v��zP�#̞|�F%d!g�6z����p�����g�B�'�z��b��B,����\�%�3��h�p/o4��a4��	:��L{|��܌��^y�V>L����JpM�R�dx��m�w���i�?�il����Ѧ���&����A��d(� ����v�a^�J�5Fq��o����h�΋SU��J�Eeȼ��{B�/�R1zS1�(-��p�<>qAO<-Z�yI�\������3+�惖ݼ�c�~���X�j�����>Ae��#O��MVg�^�r�g7j&�I>���ew+�dR@E��LKf�����1p՝Z�`v�\�ɼI8�Y-ޣ�_q'U����y������%�����	�d�%��e�0���N4Bn����ޙ3�:"�h\��J%�*�g&�B�2�� N���>�I�vm�xF��W���U��|�V��ӫ�G��֮��G?o�e�"#�s|nG4��
�KQ�$k4�<�F�T(��u�M���ߟ�BtgRӑb��7N��C&(w��8UR�����FTbG��?R�{P�}��sve�E�0c��%QX�Q1��S�{�T�o^M�����Ve0�����qDxW��ApUP�-�qo�ƓrG��	I5E��-<r�-�CN >�[�}��=ũ������8NP�hg��\n��=5g9H��Y8?��_��	�Ν^T�=��2����c�vpELG����.�����˿�W��9S7d sRu�-��j4?r���A�A�(���@HjY�7g����u�u|�d=(}ا���{f1dw=�2eMV�1J��N�ب�/*�i����2h��$�.�s66A�x�MP��.y�=�`�j����#QEZ��r�s	3����B������S�d������k�yS�{2Eq������Ty�L{�.Ć|÷M��~w��OlG6�z<#}�߷d��n4�>Z����B0K`Q�l�_���)s��=XcOi��I_�n�1�@ /E���؍��~���{8��sd�U�Su�˒~��K*�j}��u�XJ��ʷ�r*�����*���aW��D���w196�}��c�8�k����\��*�c�{|�m�''���3��]�ؚAݻ������R��A'�v�T��\�f���Ǚ�����uX����)�D,G0<7_n�_�Kv�D�� ����g��O��j��s3D���}��-0�o����E�w�O�7�.o�ӺJ;��B-k7H�+����.H=���3^��?N.����[W��������ZG-�<�. ܃�ɳ[�Q���Gi"���H+U#�c���	|�5���r*|��� ��P�F�������2@ܘm�"J���G�=�������<�v�鿊���jɀ�4rנ�`������Jv�gx����"7�h5�
�%��O��:���ZK-���ZT菔�m��D���`�+�PJ�����ӳQ�XS�������f�U���L�ͥ�F���=�@C1�IȦ��?a��J(,_="�?7;�~do�k���i+u#@+��O�? �
��p�1�J�M}e�޻a�)<5�{���Շ��vl�O�ìs�pO�����.K*����d_��s
��L���_�K�_oa{�e��:��tJ��3B�k�TyP��̵z�X������$�m�2sp�z*剣�'�Hț��g����\PFKݴ���C�Gb�VI١|����F�h��q��H�̭J��g��?h�V#��=ŉ<y��`b�罏�lys��3$ף����?7�*�M�����X��sT����(��2m�=��&��X���{4���R஬z�N��3Q�C1zR).���~���V�q }O��\�̐��*׺��;�G/B����i��*�st$�M�s��^�1�?ݻ��U�?�������lO��QU'���䕪�]�
j��=�0fuG�O�x�"�arDY����V_iܖ�5(���v	y�B�����Jݞ����[8:O~�  �l��=h�^u?���l0�̉&vW�D�w��7q"LJ�K���Ab-��Mgri+�?�Q�A[�����h�I��7i�I	��5�ԉ$�l�/��u��!�3-�shVt�ww�qOU?^��I��u��7�6��cU+���<���{�A֘U��Y�N�?PC�\��@�>�?�;�a.�ʪ�"'�!���x���H?���v�$@�|-��.+�m-	�����x��o�g�8�fz���YyoG*A���\�Qt
2]�Оk�%��Z��F��]{u���-��TTD|W��c�(�!��VpJDB�ZN3[��RZ�,��²�C�4��{���R�L.� ^ќm�G�(���JG���F��#��H��p��6�g�,5<a���8&ĀM�	���m��'�=�0�*��u_ *0i>|����g��z�I￙��S��0D��>Ct8y�K�,��e�Ѝ.��D�6#�8�v��w�C�!�Ġ��]���Av	\դ �Nh�O���((H����9���j}�a��۪T�k=��/���7��ϻ�p�yow�eCteY��/~l� � #u}�b�xdc�!���J���S,�~�j�3���\2Wn��v�v�

D(�s�ˌ������P / �@����$�!�Bt:i]�y��?��Gpdث6�Le/J���G={��ۏnxX���U@Qٰ/����^��B��v/qu���	�~� ��C�_�U��T�^'*�7N~<���Z�iS�h���܇cjg����R���2��������RnX<�f4Lғ�H�sQ-��Պ�7��t9����}�Z�I!�ݗ� D$͓��w��d@��h��9I�jB����r]r�f��()ak���OB�C�s�{�a�=����*�v*�.�hD�V��<�dpP�R��:�c�$(�߇R.�{i�KJ�P���·����v�kC�mÏ���M�퇐�g���j{be�(�����w��)�O������ �
Y��7��f��5�Aa~�e:ve��y+���3Wq*�3�����'6����q��b� '�al �S4k���UQ��y=w��!���n���jX����UXvB /멤��V�S	j���=�!ı��i�����c�R�.0Knd��ޏ�P�R9�h_K���}|T+5��R则,����BAi����F -�r�ᙊ15�۠�󬤏ld�����7�.�ѩmYN7�-��3w(�9�9so��y1��c��/i��Ƀ����.�<� �$������x8R��Y?�|��(�/p˔%�R�PLT�g�Q!�B80#v�����CE��O����VFLN�z鰍������y�0�E��b}��n4�w�Cտ�|��6�״�쨶� ���`�2�@*�a�y[,m�2J��zъ|t�]b;[`QOE+��Ko�#��I��c}F84��wS˸2��NzZ ˊ�� ���*�0�bD8Q~����f=�X����̓�UX�T�Z�V+��uem�Z���Jp�*�Ł]��g�M@ę��4��5٭2���oPݬF�' B�e�Ç�i��m0��Q"��!���1d6n�Ξ�"�����E[��%Y�V���%�����T����@B�U�����=C��i����H���a9�
l�BD�M戜�Ca�����~��X���^��@OU"�iy�����l<
Qè��1���us�*��b�!��:MA�
m��$���y��RԴ[���
A�$�a�?��{���p�>�L�.��C;No��Q�\-q�iZE�J�Y����{�:�^���O�������ju�#�|��y���������� 'j5PJ�����l/=4=��C�,ʼ��4V�&����R�E�������!�y
te��Ȗ�*�&$����$�L�oo
@�eU�-'})s\���m?� v��|S�Pܛ��۩1Z���>U�-��A����xH�Vћx5n||[�#	zuu�-�9R�Ȥ���)yF�y��B&�[��$���X�brX���-=����6![u�u�,��Q��r(�g?{�:�4+�|Ȏ�f=N9�Oe]̂�\=y�]��|8������1�́�����~���D�q6S��2[�݀��m*�r���	�r-8����F�c����������$a������ep��!��i��
w�Đ-�Hi��{-�A��HV��Q�^��K�N뼫<E�&��Tf?��z�+D�m&����l�d�K*%�N�&�5&u���b�W�����)�X4!��<��O8\(K����;�3���-�
t�&��Jv��JelZo��Ӹ!�?7�N�鯞A!tT���G�@��YE��+������x�E�5q����g�t;|)j��E[���ǐk��F)o{I�w�;4�?�%�PQp�����w�����4y<�<�3����iC��܁Ǖu/C��JW�U���g�Z��U�^�#);��lO�3O�w��Wz�����\&D���d<{�#� 8X�������Y��[r���x�t�y''��V|T�i\���-p���$�Ğy��
��V�����X�>b2´��Az%@!�<j��V�_�����n��	��\`�6�o�p[��/s?���$�g�}.��kH�GW�a�`�'D�KY����e������ i�VG�b���q���X��4��1��g�����L��8��O���Y��w��m�j�Ӯ����C�%;�1�%m���R�ZY��U��َ���Ͽ�l���})�l�����VXJ�����"D���>��*�7;����2��q���c��*���|:��|�ek)�7�nЛ�	�{���C���t��0�2Mu�����.�E듗��DWz,�z`�Ʋr�O�*��Yh]�����~���u宫 0��v�1�\�Æ*����l���-�l2�$��̚O0D�|G���=P�
B$V�>��䶏Iuvy݌�W�.[����@v��ZQ"���h�ڥ��1�w!5A{�j=��`�
Ů��S��6}�XС�y�9����پn������m�Bjݼ������X�Τ��PD}�WT��e�" fS#�wwʱ�6�J����e�:��h�#�`��9�'!
ü�<q��}�>:�2tC��d�H�V5�R�N&�]8����'��"nd�����t���ݭ2ܡ�9����=�\N�=��*�zzs* �]���y��Ņ�t�r[�82���2^-I�u��Г��E���Ch���y(������P�w���V4	����G gnJ}���޹l�e�������D,�tӱ�3y�at�xH�V���#O�p�D�Pג,�}�'^�X:�m5=��G0Q���x{Z��\ ��J��ݍ�(�����x#2W�q�ş�	��*M�mN �}�j�{V�M	i���b,k�"c�K����~v:�آE�Co���A��Oc�ZJ^s���eJ՝{�X���H�EU_II\>">zȎ�C��pZ� .��}�R�i
�e�4ݴ��L-`��yҌg W2xN�	}	��W���j=;4Po<R�����C��f���6�.���L��v�R�qs�]��SqldH��N(L��|۔��>3�����T��럣E�O` �K�ߙ�q�
�ܻ����y�G���ؼo�&�tq����E��u�`~�22�u��R&��(u�$}a��a	p���U�W
Ϛ�m�����"��'2x&��5�=���P�s�TAR���O�yy�-m�CZ��Sc~a�n�>4�$+�#�a��xՏɛ����D힉��4y����j���w�jP,��ǐ�X�;������Y��Ho炑��l���T�H�'�рFG�.�PY�Z���`�yH/���#��@��+�:��-��V�ϗ�	�ީ�(�܉6���q�*X2��x]/������UkKc���)p7,�痩D���M� NW0s�ة��4~r�����\1�R���.���K�Խ�$h�T;�͡z��dȯ� ��K�xlh� �g��������d�쾰(�v�{���GQ�_��k����ڊ*��ܼ}Nʢ���X\<H�.�Fr*m)�)��i6[@( ��H�6z]�����烕;a�ډ����3�K�������ˈ-b�{H�F#���mD��H4�c��1B�(��8R�}bQ\��(�RI^9�,/9�gU���.�ue�gO@Ý���_�2�ȥ�B���HS��gs>�	�㋢�+'-B,:6��� ]cQ��;