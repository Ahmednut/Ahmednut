XlxV64EB    15ba     850�6ghS؂�O�+�	���)@5W�s��hQ�[��p/L�������DU�̅���
��vS��2M���M(?��F;�	���������a�(���k�����F�@�YJ'ӝR��4<���؎�K�T�B��s7�d�U�-Ѐ�������`x_��)8*���+��vB9���p�+���R�8�����`5@o�`��8�h��y�*«8i�[nr+I���H���1y�u���ؠg�<�:���">�1+��SU5�]�!v]�'���$�Ew���\y�|�Ez�w��̤� Yl3�)��~��|Cf�XD��aAo�~^	���t,�x �N�����'��%��l1F�.1=��֏+2����r�Og�-r�E`�HX�"C�%2�́-�1K~�kz��1���"�Y�(Ά�{t�� ӈ� >����b��@bH$��~hUkҨ`h�Hğ+��!p\E�)쿢�6߼ueaDubt��E?P�����$$�_�iKUͰ+�t��xz٧�O�M���'�AI��w�&�9�SG)- }w�:O�w⭉\�GL>h�=��F+�ENx�o��=:�uJ�8�����ah�{�>t����H�<h��'"hm��o���k�[N�N�>�wh��Y6*�_#���v�_v��cΏ�V��_�������X�X+hY;N�	���/�=!w�;v���/É��/2_�f>	�=�e���{8�����^��^���5���gm�Tj
�jFo"/db�bt�7���.��i���'���} �[�D�[�O�䂫��~
i�BiCF]��ͥor���Ӗ�գ� ��C�~�Ҭ������$�j��F�$�`Z�c��W�kvD�Up`�&�&1�#�yxI��j��0.Թ�"��W�EF��kG|ڇ��a�ڇ)I���`18qt�",��ޕy}&
�/��>�)FY�����m���t�<��b`!���ۗ*���ISl�bbh�]2&"���xY:��O�)���@�'E�J ��ؕ�Zr�s�럥j�j��5�����������1�Fq ��Z����<]d`�Ak�����g]��M����\��h��VpƉj6��:F�Q�����`�����e� � �E�����մ���GK�
�4�����G�-���Z���=ew�-]���oK:CS�l7���w����HX��l�ߝTz�h�>�1 ����#����
=�GV�W=���G���C�����;��Gbi���&�����j��*��Zcɗ[C��F�5�{��	?EK�Ib���hi\�@	�뗠4r�"���@h��s`^��ԴV�[�������Y�X5w�=B�;��ƀ�Jh��.�׷+׻S�|��-�k`*�f߷��~��#�����$��e���Q`k6�Y���x
��1e��~أJ>��"�T���/$/���6�	�Ƣ�pC�R*L�T���[5K��ˑ������1�ɰB�x�}�44��� >�cX5��B��8�sI3���	>���UK6�t��O��ϙ6���$����譥��3X�G��+G�J��q�m�ݧ�G�	Z����%���q��r5�����2�{�<*������JI�^O6ӆ�;��G�N ��v����� �fY)m�N�k�n#�G��l$�q��󉮏����_�-��#��x����5��5Xd�io�r]Ҳ^���3}�ڥP�;a��=���h��U����=�ZG*�HTv*a�ZQ�׀tWi����0���_���lvuAR���:���<p��ڥ^oʉ,QM��
o?��I�'.\K'C�Mv������!3A4�C�h����{��h��+Џr��f�����F��-|?��h/θ�3g�b終��u*�x+\��kk��"U	�ٲ��R�r��u6�tQ�%�Qq���l�nju�K"�T��;���"M1sJb�U�l�1�gwTb�����\#/�Ll��������N��SxQ�m'["m�L����� X�;j!T���_G�4	Z��Od�P|������ }�t|l.�k�K�_#9�HгP��Lm_j��'���)���<t�