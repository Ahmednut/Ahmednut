XlxV64EB    25d9     aa0.T���缭t�#DN5NH��Da{�g���w,UA�[����"g��Q&[Z pS�mZ�#�����3w
d�y��8��{ Z@@�^"�7L�v�p|�I�T:fS�y<>�`������1���8_V�LvF�!sm����z�C}jJg���i4,�B�q��jJ��B����¹x�{����UJ�A��s�|��<�=����$XI)���-1��?6��-{Jg}6�M?�����܇[�ˏM�����OlJ��x_�X#bة�3����=�����2$�� �Q�DZ�X����	+��RaY��{�������.m�q!��F�}~�w�1�|�����R�R��A�A���T5��ձ4�Z�;�kxН�����[9�E�9sH��������sov��z{���8�S�4:4Qgi��c�q�b���<,��==�A���dŒ��&�<��p����w <ьȠ+a��d�
@b_�V͆Ĵ���K5�-�QՈ>�.�V/��ɼJ���kW�z��q�oB�����뽸fܞ�F����X�h��E��0�b��I�����ת�h����m{xr�hG͔P�@*&�������)Ex��"��ظp�0�U����Ji��Q=k���D~�w6r�pX
���gk�?�o���0�� 3)�:�3Q�� eP�\ؔ��f]����D��*�5����3�O�߰hA�ރ��P����Ezvd��f��e��wi*}a�)? �
��~*�K��cEhޤ�^-ɨ��=�t"�D�g�j�y����8m��@/E��*v5,�v��hw��F���F�1�8Q���0/a��p��fg}��o"�]n�t�)H#�GG�X��<hd�U6�z&ia.�u��㉷d0X������7i�����	
���9� U�s��^Ǝ�l�8;�هƽ��v��׳|���l1Ŷ^�"1|��r��H� �\�M�n|��]��Ȑ����?Z2�~�"�q�e��:�L!���ܟ��V:0��_��Cdٞ2*�ah�9�����t�����2��kO�8ܾ/Ow�:��[|�P���)1�Z����\���8'��8k[�֌��uX.{�?�������<�>��>tC�@+��<-�wPB���������Zq����=}�m\����^y�j��0��;�t�G�J����؏@}�k�:�,��7/�&"���n��=#�)'.�3*��ݡ֊�Ys�Te��f}Ӆ���P�oZ���n;۳�X
����}����]1��U-�.h�0[}M4)�e%�����CA��`.�@s]�%�ԉ[p]?�$Eΐ��Ȗ�[H>u�U	Hg�:�S��~80	�8|�O��cZ��Pډ8v�lќ�S�?���2�@�<��	��Vq�E�R��:��5�ې��Ɩ9i��&��������,ӆ�п�N9 
�rL��s�7.�a��U��$]^�13]�"�bق�DBk�:�E�XE#"S^�FP<EJ��ֽqc���o�Y�<�,9��t�|'���T{��Y'Q���r����¨q9��n߁*k�:�K�Ħx6ָ��9SL�I�a��Z���P���5s� i鰬�b��k�'�I����(H�r9-o���X1	#Jk/�����'q�O@lftg���}�p�� ���O�2��*�?8�Lcu9�P�TRY+CMW�~f�	#�Np�׶q$����i݌yPH!�:e�?��ѽĮ�9߱W X�R��'�_�3GK]��%65���s7�a��b���I7u/ǟ�)[�i:�}P�w̄��±�ZDQ�*�ƹ��_���J�.�%��j(��Rg�����Ƹ[�o�Xp�:�/B�Ð֕IFԭ��RM�������0�X@\f\�g2���}��Ui�b����e�LOj�Տ��Wq08����M���k�t$)�Np?������7=�_i[�k�Z7��﮺�8�f?Ha��IF:�>��)�7�Y4���	k���P7��O�r
>��`�����9�l�p��d�E�d;���OEv���q+iC�`�IW�0S�V(ʑgzJ@�s�0�e���^�`��B���4�P�9�B�@ﯸ����9K�<ޓ���� �jΪ��f��2 ��]����}t���3&kƙJ����C���ƈH�?�E�d���LD�pc{`�OI^ˍ���Q5&��駀ca�v�T�e�X|�Jn��c6>w�w����7�$��X[�)�^��|x�G��r5�3�+́,Ppԣ7	\��+����U�F�UwZ|�O��]@�q~��U�!3��w�i_7(.<�IB����1�A=z��/A=��+�� ��v���*9>oq���eRy�ٹ�8��J��=z��閦��*j�O��l�9�h��1��i����4�v�z����֯�G�����ɪW�3|8�R�"�������S�<�y�ؼ��e!�����i�i`�r�,0΀��dUc�7�J�x�%��R9�G3�"��|�b�)FB�r%g�9w����ǹ���&���o�Vʫd��oRYΞ��m$	�;�dK����l��^)�>�T*�z�4-
|.C�}2D��S@̆�Z� B���`}��یaԓ���"=�@�$���
gSêr�V�K�˪K1�;��1�K�T%�A:m	�_�� �$e4P���ha�i`��~:%�+'�}}��9�2Z�F�m�t,S���z�ȳ��%V