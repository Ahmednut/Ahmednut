--------------------------------------------------------------------------------   
-- 
--    ****                              *                                     
--   ******                            ***                                    
--   *******                           ****                                   
--   ********    ****  ****     **** *********    ******* ****    *********** 
--   *********   ****  ****     **** *********  **************  ************* 
--   **** *****  ****  ****     ****   ****    *****    ****** *****     **** 
--   ****  ***** ****  ****     ****   ****   *****      ****  ****      **** 
--  ****    *********  ****     ****   ****   ****       ****  ****      **** 
--  ****     ********  ****    *****  ****    *****     *****  ****      **** 
--  ****      ******   ***** ******   *****    ****** *******  ****** ******* 
--  ****        ****   ************    ******   *************   ************* 
--  ****         ***     ****  ****     ****      *****  ****     *****  **** 
--                                                                       **** 
--          I N N O V A T I O N  T O D A Y  F O R  T O M M O R O W       **** 
--                                                                        ***       
-- 
--------------------------------------------------------------------------------
-- Filename:          user_logic.vhd
-- Version:           v1_00_a
-- Description:       User Logic implementation module
-- Generated by:      julien.roy
-- Date:              2013-08-01 16:18:09
-- Generated:         using LyrtechRD REGGENUTIL based on Xilinx IPIF Wizard.
-- VHDL Standard:     VHDL'93
------------------------------------------------------------------------------
-- Copyright (c) 2001-2012 LYRtech RD Inc.  All rights reserved.
------------------------------------------------------------------------------
--
-----------------------------------------------------------------------------
-- Register Memory Map & Description
-----------------------------------------------------------------------------
-- BASEADDR + 0x0   MI125INFO    bits to get the MI125 info
--   15:0 Version R
--   31:16 CoreID R

-- BASEADDR + 0x4   MI125CTRL    bits to control the MI125 Inner logic
--   0:0 UpdateADCStatus P O=o_UpdateADCStatus_p
--   1:1 IdelayRst R W O=o_IdelayRst_p
--   14:10 TriggerDelay R W O=ov5_TriggerDelay_p
--   15:15 reset_calib_detection R W O=o_reset_calib_detection_p
--   2:2 IdelayCtrlRst R W O=o_IdelayCtrlRst_p
--   3:3 IserdesRst R W O=o_IserdesRst_p
--   31:16 AdcValid R W O=ov16_AdcValid_p
--   4:4 DigOutRandEn R W O=o_DigOutRandEn_p
--   5:5 IPSoftRst R W O=o_IPSoftRst_p
--   7:6 ChannelConfig R W O=ov2_ChannelConfig_p
--   8:8 DataFormat R W O=o_DataFormat_p
--   9:9 ADCClockMMCMRst R W O=o_ADCClockMMCMRst_p

-- BASEADDR + 0x8   MI125STATUS    General status register
--   0:0 idelay_ready R I=i_idelay_ready_p
--   1:1 calib_detection_done R I=i_calib_detection_done_p
--   2:2 ADCClockMMCMLocked R I=i_ADCClockMMCMLocked_p
--   3:3 ADCClockMMCMPresent R I=i_ADCClockMMCMPresent_p
--   31:8 rsvd2 R
--   7:4 FmcPosition R I=iv4_FmcPosition_p

-- BASEADDR + 0xc   MI125ADCIDELAYVALUE    adc Idelay Value
--   31:10 rsvd R
--   4:0 adcIdelay_value R W O=ov5_adcIdelay_value_p
--   9:5 clkIdelay_value R W O=ov5_clkIdelay_value_p

-- BASEADDR + 0x10   MI125ADCIDELAYWE   adc Idelay mask
--   31:0 adcIdelay_we P O=ov32_adcIdelay_we_p

-- BASEADDR + 0x14   MI125BITSLIP   bitslip mask
--   31:0 bitslip P O=ov32_bitslip_p

-- BASEADDR + 0x18   MI125CALIBERROR   Indicate if the data is stable for each lane
--   31:0 calib_error R I=iv32_calib_error_p

-- BASEADDR + 0x1c   MI125CALIBPATTERNERROR   Indicate if the data is the same than the calibration pattern for each lane
--   31:0 calib_pattern_error R I=iv32_calib_pattern_error_p

-- BASEADDR + 0x20   MI125FREQCNTCLK   Control and status of the clock frequency counter
--   15:0 FreqCntClkCnt R I=iv16_FreqCntClkCnt_p
--   21:16 FreqCntClkSel R W O=ov6_FreqCntClkSel_p
--   22:22 FreqCntRst R W O=o_FreqCntRst_p
--   31:23 rsvd R

--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library proc_common_v3_00_a;
use proc_common_v3_00_a.proc_common_pkg.all;

-- DO NOT EDIT ABOVE THIS LINE --------------------

--USER libraries added here

------------------------------------------------------------------------------
-- Entity section
------------------------------------------------------------------------------
-- Definition of Generics:
--   C_NUM_REG                    -- Number of software accessible registers
--   C_SLV_DWIDTH                 -- Slave interface data bus width
--
-- Definition of Ports:
--   Bus2IP_Clk                   -- Bus to IP clock
--   Bus2IP_Resetn                -- Bus to IP reset
--   Bus2IP_Data                  -- Bus to IP data bus
--   Bus2IP_BE                    -- Bus to IP byte enables
--   Bus2IP_RdCE                  -- Bus to IP read chip enable
--   Bus2IP_WrCE                  -- Bus to IP write chip enable
--   IP2Bus_Data                  -- IP to Bus data bus
--   IP2Bus_RdAck                 -- IP to Bus read transfer acknowledgement
--   IP2Bus_WrAck                 -- IP to Bus write transfer acknowledgement
--   IP2Bus_Error                 -- IP to Bus error response
------------------------------------------------------------------------------

entity user_logic is
  generic
  (
    -- ADD USER GENERICS BELOW THIS LINE ---------------
    --USER generics added here
    -- ADD USER GENERICS ABOVE THIS LINE ---------------
    C_BUILD_REVISION               : std_logic_vector := X"0000";
    -- DO NOT EDIT BELOW THIS LINE ---------------------
    -- Bus protocol parameters, do not add to or delete
    C_NUM_REG                      : integer              := 9;
    C_SLV_DWIDTH                   : integer              := 32
    -- DO NOT EDIT ABOVE THIS LINE ---------------------
  );
  port
  (
    -- ADD USER PORTS BELOW THIS LINE ------------------
    --USER ports added here
    -- ADD USER PORTS ABOVE THIS LINE ------------------
    -- User ports
    i_logicRst_p : in std_logic;

    o_UpdateADCStatus_p : out std_logic;
    o_IdelayRst_p : out std_logic;
    ov5_TriggerDelay_p : out std_logic_vector(4 downto 0);
    o_reset_calib_detection_p : out std_logic;
    o_IdelayCtrlRst_p : out std_logic;
    o_IserdesRst_p : out std_logic;
    ov16_AdcValid_p : out std_logic_vector(15 downto 0);
    o_DigOutRandEn_p : out std_logic;
    o_IPSoftRst_p : out std_logic;
    ov2_ChannelConfig_p : out std_logic_vector(1 downto 0);
    o_DataFormat_p : out std_logic;
    o_ADCClockMMCMRst_p : out std_logic;
    i_idelay_ready_p : in std_logic;
    i_calib_detection_done_p : in std_logic;
    i_ADCClockMMCMLocked_p : in std_logic;
    i_ADCClockMMCMPresent_p : in std_logic;
    iv4_FmcPosition_p : in std_logic_vector(3 downto 0);
    ov5_adcIdelay_value_p : out std_logic_vector(4 downto 0);
    ov5_clkIdelay_value_p : out std_logic_vector(4 downto 0);
    ov32_adcIdelay_we_p : out std_logic_vector(31 downto 0);
    ov32_bitslip_p : out std_logic_vector(31 downto 0);
    iv32_calib_error_p : in std_logic_vector(31 downto 0);
    iv32_calib_pattern_error_p : in std_logic_vector(31 downto 0);
    iv16_FreqCntClkCnt_p : in std_logic_vector(15 downto 0);
    ov6_FreqCntClkSel_p : out std_logic_vector(5 downto 0);
    o_FreqCntRst_p : out std_logic;
    -- Bus protocol ports, do not add to or delete
    Bus2IP_Clk                     : in  std_logic;
    Bus2IP_Resetn                  : in  std_logic;
    Bus2IP_Data                    : in  std_logic_vector(C_SLV_DWIDTH-1 downto 0);
    Bus2IP_BE                      : in  std_logic_vector(C_SLV_DWIDTH/8-1 downto 0);
    Bus2IP_RdCE                    : in  std_logic_vector(C_NUM_REG-1 downto 0);
    Bus2IP_WrCE                    : in  std_logic_vector(C_NUM_REG-1 downto 0);
    IP2Bus_Data                    : out std_logic_vector(C_SLV_DWIDTH-1 downto 0);
    IP2Bus_RdAck                   : out std_logic;
    IP2Bus_WrAck                   : out std_logic;
    IP2Bus_Error                   : out std_logic
  );

 attribute MAX_FANOUT : string;
 attribute SIGIS : string;
 attribute SIGIS of Bus2IP_Clk    : signal is "CLK";
 attribute SIGIS of Bus2IP_Resetn : signal is "RST";

end entity user_logic;

------------------------------------------------------------------------------
-- Architecture section
------------------------------------------------------------------------------

architecture IMP of user_logic is

-------------------------------------------------------------------------------
-- Constant declarations
-------------------------------------------------------------------------------


-------------------------------------------------------------------------------
--     ************** Function declaratin *******************                   
-- Return a std_logic_vector with only one bit set to one.
-- The argument BitPosition represent the bit position to set to one, starting with 0.
-- The argument Width represent the width of the returned std_logic_vector.
-------------------------------------------------------------------------------
  function OneHotVector( BitPosition : integer;                              
                Width : integer)                                             
                return std_logic_vector                                      
  is                                                                         
    variable Result                   : std_logic_vector(Width - 1 downto 0);

  begin                        
    Result := (others => '0'); 
    Result(BitPosition) := '1';
    return Result;             
  end OneHotVector;            
-------------------------------------------------------------------------------
-- Signal and Type Declarations
-------------------------------------------------------------------------------

  signal UpdateADCStatus_s                     : std_logic;
  signal IdelayRst_s                     : std_logic;
  signal v5_TriggerDelay_s                     : std_logic_vector(4 downto 0);
  signal reset_calib_detection_s                     : std_logic;
  signal IdelayCtrlRst_s                     : std_logic;
  signal IserdesRst_s                     : std_logic;
  signal v16_AdcValid_s                     : std_logic_vector(15 downto 0);
  signal DigOutRandEn_s                     : std_logic;
  signal IPSoftRst_s                     : std_logic;
  signal v2_ChannelConfig_s                     : std_logic_vector(1 downto 0);
  signal DataFormat_s                     : std_logic;
  signal ADCClockMMCMRst_s                     : std_logic;
  signal v5_adcIdelay_value_s                     : std_logic_vector(4 downto 0);
  signal v5_clkIdelay_value_s                     : std_logic_vector(4 downto 0);
  signal v32_adcIdelay_we_s                     : std_logic_vector(31 downto 0);
  signal v32_bitslip_s                     : std_logic_vector(31 downto 0);
  signal v6_FreqCntClkSel_s                     : std_logic_vector(5 downto 0);
  signal FreqCntRst_s                     : std_logic;
  signal slv_reg_write_sel              : std_logic_vector(8 downto 0);
  signal slv_reg_read_sel               : std_logic_vector(8 downto 0);
  signal slv_ip2bus_data                : std_logic_vector(C_SLV_DWIDTH-1 downto 0);
  signal slv_read_ack                   : std_logic;
  signal slv_write_ack                  : std_logic;
  
  attribute KEEP : string;
  attribute KEEP of IPSoftRst_s : signal is "TRUE";    

------------------------------------------------------------------------------
begin
------------------------------------------------------------------------------

-------------------------------------------------------------------------------
-- Begin architecture
-------------------------------------------------------------------------------

-- swap bits
WrCeBitSwap: for i in 0 to slv_reg_write_sel'high generate
  slv_reg_write_sel(i) <= Bus2IP_WrCE(slv_reg_write_sel'high - i);
end generate WrCeBitSwap;

RdCeBitSwap: for i in 0 to slv_reg_read_sel'high generate
  slv_reg_read_sel(i)  <= Bus2IP_RdCE(slv_reg_read_sel'high - i);
end generate RdCeBitSwap;

-- generate write/read ack
  slv_write_ack <=   Bus2IP_WrCE(0) or   Bus2IP_WrCE(1) or   Bus2IP_WrCE(2) or   Bus2IP_WrCE(3) or   Bus2IP_WrCE(4) or   Bus2IP_WrCE(5) or   Bus2IP_WrCE(6) or   Bus2IP_WrCE(7) or   Bus2IP_WrCE(8);
  slv_read_ack  <=   Bus2IP_RdCE(0) or   Bus2IP_RdCE(1) or   Bus2IP_RdCE(2) or   Bus2IP_RdCE(3) or   Bus2IP_RdCE(4) or   Bus2IP_RdCE(5) or   Bus2IP_RdCE(6) or   Bus2IP_RdCE(7) or   Bus2IP_RdCE(8);

 -- implement slave model software accessible register(s)
 SLAVE_REG_WRITE_PROC : process( Bus2IP_Clk ) is
 begin

  if Bus2IP_Clk'event and Bus2IP_Clk = '1' then
    if Bus2IP_Resetn = '0' then
      UpdateADCStatus_s <= '0';
      IdelayRst_s <= '1';
      v5_TriggerDelay_s <= "00111";
      reset_calib_detection_s <= '1';
      IdelayCtrlRst_s <= '1';
      IserdesRst_s <= '1';
      v16_AdcValid_s <= "0000000000000000";
      DigOutRandEn_s <= '0';
      IPSoftRst_s <= '1';
      v2_ChannelConfig_s <= "11";
      DataFormat_s <= '1';
      ADCClockMMCMRst_s <= '0';
      v5_adcIdelay_value_s <= "00000";
      v5_clkIdelay_value_s <= "00000";
      v32_adcIdelay_we_s <= X"00000000";
      v32_bitslip_s <= X"00000000";
      v6_FreqCntClkSel_s <= "000000";
      FreqCntRst_s <= '0';

    else

  -- Synchronous reset
  if ( i_logicRst_p = '1' ) then
    UpdateADCStatus_s <= '0';
    IdelayRst_s <= '1';
    v5_TriggerDelay_s <= "00111";
    reset_calib_detection_s <= '1';
    IdelayCtrlRst_s <= '1';
    IserdesRst_s <= '1';
    v16_AdcValid_s <= "0000000000000000";
    DigOutRandEn_s <= '0';
    IPSoftRst_s <= '1';
    v2_ChannelConfig_s <= "11";
    DataFormat_s <= '1';
    ADCClockMMCMRst_s <= '0';
    v5_adcIdelay_value_s <= "00000";
    v5_clkIdelay_value_s <= "00000";
    v32_adcIdelay_we_s <= X"00000000";
    v32_bitslip_s <= X"00000000";
    v6_FreqCntClkSel_s <= "000000";
    FreqCntRst_s <= '0';
  end if;

  UpdateADCStatus_s <= '0';
  v32_adcIdelay_we_s <= X"00000000";
  v32_bitslip_s <= X"00000000";
      case slv_reg_write_sel is

        when OneHotVector(1,9) =>
          if (Bus2IP_BE(0) = '1') then
            UpdateADCStatus_s <= Bus2IP_Data(0);
          end if;
          if (Bus2IP_BE(0) = '1') then
            IdelayRst_s <= Bus2IP_Data(1);
          end if;
          if (Bus2IP_BE(1) = '1') then
            v5_TriggerDelay_s <= Bus2IP_Data(14 downto 10);
          end if;
          if (Bus2IP_BE(1) = '1') then
            reset_calib_detection_s <= Bus2IP_Data(15);
          end if;
          if (Bus2IP_BE(0) = '1') then
            IdelayCtrlRst_s <= Bus2IP_Data(2);
          end if;
          if (Bus2IP_BE(0) = '1') then
            IserdesRst_s <= Bus2IP_Data(3);
          end if;
          if (Bus2IP_BE(2) = '1') then
            v16_AdcValid_s(7 downto 0) <= Bus2IP_Data(23 downto 16);
          end if;
          if (Bus2IP_BE(3) = '1') then
            v16_AdcValid_s(15 downto 8) <= Bus2IP_Data(31 downto 24);
          end if;
          if (Bus2IP_BE(0) = '1') then
            DigOutRandEn_s <= Bus2IP_Data(4);
          end if;
          if (Bus2IP_BE(0) = '1') then
            IPSoftRst_s <= Bus2IP_Data(5);
          end if;
          if (Bus2IP_BE(0) = '1') then
            v2_ChannelConfig_s <= Bus2IP_Data(7 downto 6);
          end if;
          if (Bus2IP_BE(1) = '1') then
            DataFormat_s <= Bus2IP_Data(8);
          end if;
          if (Bus2IP_BE(1) = '1') then
            ADCClockMMCMRst_s <= Bus2IP_Data(9);
          end if;

        when OneHotVector(3,9) =>
          if (Bus2IP_BE(0) = '1') then
            v5_adcIdelay_value_s <= Bus2IP_Data(4 downto 0);
          end if;
          if (Bus2IP_BE(0) = '1') then
            v5_clkIdelay_value_s(2 downto 0) <= Bus2IP_Data(7 downto 5);
          end if;
          if (Bus2IP_BE(1) = '1') then
            v5_clkIdelay_value_s(4 downto 3) <= Bus2IP_Data(9 downto 8);
          end if;

        when OneHotVector(4,9) =>
          if (Bus2IP_BE(0) = '1') then
            v32_adcIdelay_we_s(7 downto 0) <= Bus2IP_Data(7 downto 0);
          end if;
          if (Bus2IP_BE(1) = '1') then
            v32_adcIdelay_we_s(15 downto 8) <= Bus2IP_Data(15 downto 8);
          end if;
          if (Bus2IP_BE(2) = '1') then
            v32_adcIdelay_we_s(23 downto 16) <= Bus2IP_Data(23 downto 16);
          end if;
          if (Bus2IP_BE(3) = '1') then
            v32_adcIdelay_we_s(31 downto 24) <= Bus2IP_Data(31 downto 24);
          end if;

        when OneHotVector(5,9) =>
          if (Bus2IP_BE(0) = '1') then
            v32_bitslip_s(7 downto 0) <= Bus2IP_Data(7 downto 0);
          end if;
          if (Bus2IP_BE(1) = '1') then
            v32_bitslip_s(15 downto 8) <= Bus2IP_Data(15 downto 8);
          end if;
          if (Bus2IP_BE(2) = '1') then
            v32_bitslip_s(23 downto 16) <= Bus2IP_Data(23 downto 16);
          end if;
          if (Bus2IP_BE(3) = '1') then
            v32_bitslip_s(31 downto 24) <= Bus2IP_Data(31 downto 24);
          end if;

        when OneHotVector(8,9) =>
          if (Bus2IP_BE(2) = '1') then
            v6_FreqCntClkSel_s <= Bus2IP_Data(21 downto 16);
          end if;
          if (Bus2IP_BE(2) = '1') then
            FreqCntRst_s <= Bus2IP_Data(22);
          end if;
        when others =>
          null;
      end case;
    end if;
  end if;

 end process SLAVE_REG_WRITE_PROC;

 -- implement slave model software accessible register(s) read mux
SLAVE_REG_READ_PROC : process( slv_reg_read_sel, IdelayRst_s, v5_TriggerDelay_s, reset_calib_detection_s, IdelayCtrlRst_s, IserdesRst_s, v16_AdcValid_s, DigOutRandEn_s, IPSoftRst_s, v2_ChannelConfig_s, DataFormat_s, ADCClockMMCMRst_s, i_idelay_ready_p, i_calib_detection_done_p, i_ADCClockMMCMLocked_p, i_ADCClockMMCMPresent_p, iv4_FmcPosition_p, v5_adcIdelay_value_s, iv32_calib_error_p, iv32_calib_pattern_error_p, iv16_FreqCntClkCnt_p, v6_FreqCntClkSel_s, FreqCntRst_s) is
 begin
   case slv_reg_read_sel is

        when OneHotVector(0,9) =>
          slv_ip2bus_data(15 downto 0) <= C_BUILD_REVISION;
          slv_ip2bus_data(31 downto 16) <= X"C125";

        when OneHotVector(1,9) =>
          slv_ip2bus_data(1) <= IdelayRst_s;
          slv_ip2bus_data(14 downto 10) <= v5_TriggerDelay_s;
          slv_ip2bus_data(15) <= reset_calib_detection_s;
          slv_ip2bus_data(2) <= IdelayCtrlRst_s;
          slv_ip2bus_data(3) <= IserdesRst_s;
          slv_ip2bus_data(31 downto 16) <= v16_AdcValid_s;
          slv_ip2bus_data(4) <= DigOutRandEn_s;
          slv_ip2bus_data(5) <= IPSoftRst_s;
          slv_ip2bus_data(7 downto 6) <= v2_ChannelConfig_s;
          slv_ip2bus_data(8) <= DataFormat_s;
          slv_ip2bus_data(9) <= ADCClockMMCMRst_s;

        when OneHotVector(2,9) =>
          slv_ip2bus_data(0) <= i_idelay_ready_p;
          slv_ip2bus_data(1) <= i_calib_detection_done_p;
          slv_ip2bus_data(2) <= i_ADCClockMMCMLocked_p;
          slv_ip2bus_data(3) <= i_ADCClockMMCMPresent_p;
          slv_ip2bus_data(31 downto 8) <= "000000000000000000000000";
          slv_ip2bus_data(7 downto 4) <= iv4_FmcPosition_p;

        when OneHotVector(3,9) =>
          slv_ip2bus_data(31 downto 10) <= "0000000000000000000000";
          slv_ip2bus_data(4 downto 0) <= v5_adcIdelay_value_s;
          slv_ip2bus_data(9 downto 5) <= v5_clkIdelay_value_s;

        when OneHotVector(6,9) =>
          slv_ip2bus_data(31 downto 0) <= iv32_calib_error_p;

        when OneHotVector(7,9) =>
          slv_ip2bus_data(31 downto 0) <= iv32_calib_pattern_error_p;

        when OneHotVector(8,9) =>
          slv_ip2bus_data(15 downto 0) <= iv16_FreqCntClkCnt_p;
          slv_ip2bus_data(21 downto 16) <= v6_FreqCntClkSel_s;
          slv_ip2bus_data(22) <= FreqCntRst_s;
          slv_ip2bus_data(31 downto 23) <= "000000000";
        when others =>
          slv_ip2bus_data <= (others => '0');
      end case;

 end process SLAVE_REG_READ_PROC;

------------------------------------------
-- drive IP to Bus signals
------------------------------------------
IP2Bus_Data  <= slv_ip2bus_data when slv_read_ack = '1' else (others => '0');
IP2Bus_WrAck <= slv_write_ack;
IP2Bus_RdAck <= slv_read_ack;
IP2Bus_Error <= '0';

------------------------------------------
-- Output assignments
------------------------------------------
o_UpdateADCStatus_p <= UpdateADCStatus_s;
o_IdelayRst_p <= IdelayRst_s;
ov5_TriggerDelay_p <= v5_TriggerDelay_s;
o_reset_calib_detection_p <= reset_calib_detection_s;
o_IdelayCtrlRst_p <= IdelayCtrlRst_s;
o_IserdesRst_p <= IserdesRst_s;
ov16_AdcValid_p <= v16_AdcValid_s;
o_DigOutRandEn_p <= DigOutRandEn_s;
o_IPSoftRst_p <= IPSoftRst_s;
ov2_ChannelConfig_p <= v2_ChannelConfig_s;
o_DataFormat_p <= DataFormat_s;
o_ADCClockMMCMRst_p <= ADCClockMMCMRst_s;
ov5_adcIdelay_value_p <= v5_adcIdelay_value_s;
ov5_clkIdelay_value_p <= v5_clkIdelay_value_s;
ov32_adcIdelay_we_p <= v32_adcIdelay_we_s;
ov32_bitslip_p <= v32_bitslip_s;
ov6_FreqCntClkSel_p <= v6_FreqCntClkSel_s;
o_FreqCntRst_p <= FreqCntRst_s;

end IMP;

