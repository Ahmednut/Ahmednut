XlxV64EB    fa00    22f0�~g),g�����lȨ<�OT�GϏ����R#5��R�������Me�9[�,����]�Mh=�W�0�C|ٷ���J�_��'m�C�0"�lc�:�����A��Ȕ[��e�ώ����!n�٣�wY&�0W9
�a�}�������\���r1��]�'��m#hu�v\���T�X��%��~I]�ly���
;t�@S�m�w�b�_������l���#7C����z�VZ�q��h'U�m���S�8
F����e+RdYikNf�bS�_�@ ��[��PA�������-�"/r$����n�b���v��t�غ��6�&�Ή
i�Rk�Y�U���r(���Ȩ�ms����+ͅƚV sH? S�z?"�6��k�7(��?��ӦFz.˯�#=�|�b����/h���e��,B��� �c<nJ��(��/$�����"���x��{3��;4޶����ގx��I&6��|�a^ `-�]��OĊ�|؟���Ȳ.�
��^P6*��gӺZ�Q���]'��g����U����[��z��Aޟ��G��Tq��|Yȶ�Xu��z��U'R�pkUCƑ�u`��8k=M><�ڬ�z�Z|Cˍ��Q���a�H1.7֩,����
�tt>�bg�1>�V^7KĜ�>��p��FQ+�C��-��#7P�s���!�Рx��r�-��|����G��z�y6Ȗ봕of�z�B �N�X��_.�j\��%k�^D,~�t�1�0�ÿKQ�rC99�d�iQx!&)r#!`0}�aL]���E^����K�oR�Nٳ_�}�d�-=����+�2c�Ɩ����C�-�`�wt�AH/�<(����X֌�G,tXYb5O��_�|����Oo1�B�G�,�X����l��+���A$�j�> Ve��X�Gy�yʜ�O���x��S��ۖ�%���j֟� ���CT����2Rؔ��\/�.�/f�sb��"��x̑D�[�D%p�B�0+NJ�?U,�៽̻�/9�����t��_�נE�Gt�tC�ZF��5{F<e�*��F2 ��x�ޏ��XE��v7m��z����[�>���2 �ĸ�=����
�px�&��P4�SH�L+u�(Âk���q��^�#A`����ń�|����2Ih������
r��.>'\g�ͯ���vn��d�-��P8l���p��s\����[�:�8BK߳Eu�^�!Y1��<ق7�W+܎���������+�_��������A!Y��f�lBr�lڢم:�@�b�z�yY�a�L�E��xv��WdV�8��0aU��۞r����nJ��/�X�y��/�~H�'�2T���&y�D��ᦋ��/���K����{� �	>Rp@��&,5|0�Á��?���|�`��~�j����1���)�U߾h^5	����	�M���90�4��_���=[R�N��A	DA6�$n�'(�)ܚ	l��uSP�ȤЊOU#x�	�
��RD�<[�/�i�-	�qf�P��pƼ�C6������*ȥ7��HdRè�~�1�r;]�)��T�;9"�h6�Rݹ�`�r��T����n>c�X-E����-B���X����g�{��	8�`�f]�l�&��|�o��i�M�(��mEr��t ����O�\��ą��?l�9��V�~�?ADۓ���W�m�c]��7砝���Ig�x�o��a��8B��]�����Y)JG��E��I��G���%�H�b΂*&�د�ְ��s�W�^�Y�Gˑ[\8�kFL��꿤�Ǩ�sB�;
L=����g�|�D�c�j�Y �`��R9f���h����]THUQ|�B�T��S�=��$�	�*p�
���؄d��)�a�-�nP{f�7���o"�s��x�kp��<���,4�5A ө��f�@1�Y�㈿X�-����J2��ӓ��Q�J=�"̟l<�8���Fɠ.����S���u����r�Q��g����,�p���o�t��ڈX-���{TՔq�J�	Z1q��v��v�\��ɋ���"N�����eZ����%/�n�?Dl���иi��{,^�_�XR�]$a�`����(Y���t`�&^"�J;��J��)!�`s\s��+	i͏E�hE�$�N*���> ���4�P=c=���>#��$H��ȗC�V*R�����YI$�566RO�� ^��̼r�o>N�sT���YӰ�.���Sj� �T*�
�k��2�!*�iN�S��Q�N�v��b>��M�E?�v�x�t�\�4=��~s�Z�orV�4�q<~��Q:�x+�}���7�j��q^��7��+�ɗ��˹��Vg!����K�Ew>Aą+�8�͊��E7#�8�>	^2�;M�0�ߡ�.��u|�V�1��F{q��~�W��A/�q*tg�����5[�27�Jޯ,fQt.�7�ڻG�C����՘�C�gd����E��71�j����Ӥ��0.$ohY��{�!&���,T=X�ĸw��n�!��''X¿OFF׆�*p[���Qe��V�*���,g�U�8I���%����sO[2$��� 0F��8��p�3���;k��Z�N��;ӓ��Ė��>�'�x�X��P���y_��I�,6�yn���E*���,ς�$� 0e#��k�wд�^$9��5�"���ګN�9�q�t/�[��׎�K J�q5�	>�ȩ={�Z���X��v�N���� j�����
�Jt���ߗ�� �f�(<M���oiO
 �n�X3� >1C9c+#��aL'bU���"�ܯk�r����?c�L�^~pO��g"*fJ@I��t!{k�����=\��V,@�+�ƌ�(\�i|U������.%&�?V���y�̅4c�yOF�q��o��V�
�}JO���x�(�?�_��I�19�9�EP`�s��{m��\޼������Y�-9앞7Pd��s!Q�>
4�LF��f�R���1$g @��f˩��fT?�P��k	HmE��1�'��9^��ӣ�l�i����^3��qȯ��)cZ@�-�9���uM�زv����m1����̖�����G��l`�=��^���f���i�-�é9P0�G�ӻ�I��1��׉l�m�I]�8��6B��H�·�F���?�TX�TK����u�����<�����L��Q���H�+�	\��L!`���ik�����c&i.�t6�lC`�+N.�v����  �J�M�,e�j(F[�Q�9�rҞ��x���ƺo�y@�+���4�e��O?Ri�+9��U�g��ͼ��U�m��� ����3����):�6~0=\���J[鶖˖=���G����܉+7P|��tO&�1=��ϙq�|��������]<
��o� �B H��tL���:�&s�ʟ2��q6=C� �S�����K�T���?�om�%F�˖sۖ�����j�򪼼��b|���ǲՙ-=脵��֢0D�d�O�0��)��/��G����v�#��-��%�6w� p���@\�[?f'�M�ã����*���`mYЂB��m���b�\��җ)l�X�J�Rh/��̦ �;�T9�
Fq�Ԃ���������Au�8)�����9�!����	�H��Uv��v�USP�闐��������6<ر.�L_E�%����U2�~'�×��a�����D
���]�5h��"N�Y"�#|p��%S��_���|ȡ:�e#"�M��OnSݥ'�N*A�zq����Gvg�%�>�y ����T/�8%W��L����P�J��\q���&m&�����r��oL��Oy�A��,�/] eyj�.��&�=O�%���>�r�����8u�ɬ����6t53�q^���b.ri���8��@oP��&��)���a�K�[�I�Q�:X�*�r�a�W��>�-��X� <g������o8�g+��������ʃ~䆱�S+�̐Xַ�=!-w���@=�� ��<qNYX���P;��M��XU�p�U�aY�7өʣ��0 9ep/N��w���{��W�a�n/Q�go���%�"8�WS'��X%�+\�.�R�d�_�؅���a�����~[��ӧ���l�2V�K4p���d�����V�$�
Y�����A���%H�9��$�YT�����j�J	�2L���Db=�uE-���\\t�\��ؐ8�NJV�5�`@���pKW`	�V)ff(��H��S@�Gݫ�5(m�)jrq�
~�����t���.�&$uW6	��s�P��#�Kf7�'�����t�/�'|i�ŃT8@���k��%��4s�V�7O,>�9� ��:%���[�%,-��uNE��m�1�E �ބr�J�Ԥ��N1e��>��7�,���# }��x�w����m-B!*���c(o�aՌ�̩�:��?
�'����X�{���+�lL�\ؤ��Ƥw��q���N�
6�=�}s��>�+>�p>|Ǻ�#,�!��O��( � bFu�K������j�q���W�3 I슺<�$�F�IFf��A�,�i+���2,�/5��-�L��lu��E�wT)4����=���m슎����?U �4D�t��Bv`���=��al�[��=72� -A���8��� 8s@�5��A}#J(�# +Q�B�ƺR�c��ˋ��z�h��P�PN*3��3�aEˎb��[>��2�1�&��n7K@�{� #p�g��BYIn�����TǒlXX~Ox�pɉ������Ñ��tIF���X9���A���A;�(�Á�8��7���	~� 7H:JPm��hQA�w�*����-�����}-�1G��cT�SҲ�C40Ye�j��͇>�N���	���< 1݅��VZ�����o%�į�u�nB���Z{1Z����޸�o����CneN,qGH���d���6q����FY�5x�,Q��S��G�w��8�x����D�c3٢�;a�Ŕq2_�@�.~~������HQ�WU���
�=��2�[s�,�D�}�P�&`��:T��?ԚJx9a��i�Aw�w_��4���=��H��T��[�+�720�-�fA������E����e~����@u�s)��%D�r���Z,5C�?X�"@ۊ@�go~��D����z;�2�6�HS�� 9�_2gZ��'�i�!ІJ��K� ��F�]��7�-N5kq"��z_ -�֢<=|�
��amGธ��x%&�X'x��AG�f�t�g�����X�p��''�ŸF��X5�8 �mc��y��;��ȄP?7(�(y�,����x�@��������.���T��G���,ۼ^m ~��lP�nY�y�h�������5t�X���TCI��̴kw�M.�\��ϔ?=�	�����mG�
B�9\�[�Q@�߂��M1��$b}���>�t���ֵhJ�أ�-�!Q��������I���G������%ԍ2��!j����3�|���K�L];H�{t�z�|�%���_��{����0��tTJ��F"Z��Z��OXeœ�I��T���R�Q&�%��[:ti.��˹�Ul�S��:���W�����p-�rʸf�!0�#~E�\ '��Nxo�a�ch��~_������Iŋ���#r�Q�T=�%#uH��m���`�����_�`�����W'/�9�C Ur*a����O������/���8ZW'u?k��<4D��{�0H�l��_V�<�I�ہ��mL/j�N��@���8;�����v�N�ۊ��?Ƹ.�A6����hcg�VU���>�#R����.Z�l�=/�%# �Dc�����,�u��˖=rv�f��~�o��$��O��3(��=e�=�&�w����a��������D~+k�&�ƹ����Q١�0�\���:óN�W�V0� ���Z�
�见�������e����k;4I��U!��9�ݽ�c���N�$��	��r�ʿ���Q�L������9X�l��4&�p̴����2$?�j8g�z<G]0[n$V*A{aH�x���T���_6��(���m�ܞU�/�i���f���m|=_?���f�"9c"�� �jk3�&J�'��$��g��pln��I���M�"�l����47mF2j���!j��s���B_�ϔ>� ������kS�h����~���S©n�1������	����^�_M��/��2���أ��w��d���Z1(Q���N�����ǫ���������$���F}��K�Z�E�s��2�O��m�c	��A������Kaw��^&g��A���Aĵ�aY�v��e!آŊ�ǒ�W�)K:ޞ� �H��v�诼}�����H����;n�[��r��z��$va�JId��� x�R9��3[���`agy���!�w�2wuG^YC��;KIk��oH4�>ƞ�{�+n���&9�
��Έ
yg���JK�_�~�9+�%w��)�l\A����*�x{L�S[�mR���m���~B�$h[����~�~�b"TN�|X��I�e`�g�|;ep!���E�����9,!����'�\�%��x���QD\_ڎl��Bf���=���������,���z%��rb��V���g�ގP!}ү���j����Ë1U?�E븕?�⡴�fՌ�u��nNw�����p���h|ȕ������k-6O��_���?����J4���)�ś<���+�iU��\�ݟq<�C�tX��o㨢5�[��X��&p/��OM�m���w�/r \ݣ�D�9�զH����HB���O�z������$G�,��+n���Ms�d.����>��[v�fi���-%v������Q�	���&���M��8-s9i����n�
��OC�iP�7VjE=R����#[y��,tF���?)I��X�YHAWav<�o,�_"������N�6`��xϐ�֚����$pQMe@�+_:[���ɍ�[�ݔ]�8��uK)��r�Q��v�6�j�/���D���6���n�j z����J��R���}T̖<�W�?�{�{߽�qFDn5V*�=��5W�q �U`��4v\3�.�G�Ƽh�&�w��;��Y���N�j���ފ&��]0�ֱ#D�7���0M�u��z��*7Yk ̸�ۨ{���C���W�G3�'�j%��p����f�)�|��إ(�:�������:�D�:;m�Oˀ�z�����������,Y�h�(�i���^��ۢ��(!�j$�Ċ�����޵yeII�%[�M���Y�6X
�PQ�;����#R�:UP9%���X!5Aq؜8}��F�[�����wf�[��g
�.�A�����66��停��R��K,� ��-	K����u{X��25����k�|��X�������So��|��+���9R<�M/�4�=ϳ�ACӮ��FY���-�]M5��y�>����/���Q�{<Ʉ��9Y��u��^�o/ʴ�#�ev�-��l�I��6��b�H���:.s:)��>1�cF���\������k25�)d�%?�4ށI\@�gv*�K�ﮊm���Yh��4LJa�������]o��]dh�" Z��4/�x!��Ԅ0s�#7�(����c���O͉t&O�3��7;�V���z|��D����Q&ST!��Ӿ�#����s�1s
���0H U���2�z�v�?��P���
��<B��5J
�~{��sS���o�q�L��_��f�n)�P|�-�����1n�Y��%^���[%h~}� 䲚���ɛ������y����1�������X�-;y����d=A��ug���xO�3�l�_��lћ7AM�;nX��Vi�o
�F����r�hz&�^�����'�A�:����$l��EF>�
:~OT��^"���� p8�C#Qq<B�Js(�n�H�y��N�6G<�n�%�M?�?��Yڬ�萝6�HO�ɐ'��I����'y;����q��_�!r�ׄ���iYQC�s�d'��$Ȍ&"m:3y�k�'��GfABd����A����x_L���|hw��6��'��:��φ:����2w�~-lyp�s��ɿ�K�zZkLq�6�%1�f�H��y^
�b�"8J���T�� }1!M��3a�uu�z��y  IB�_����2ת�	�\"�7�`�	�q�('M�p����*�G@����߰��)8��͙��w���Z��e��DF�c#Q���z�5������2�h~bE���V��LC8���m�E�O�f��� >Q{g Q���M�f)��	x�S���+~���KI� �ؾm	�!\� h0U@�>�W��Tۙ��� �� �~�֋Xi`���}ߢ�Xj7��0�mf��|���7좤ø�\�F=��,�J�`��X�A'��Ĺ��������ck�%D�XAo��dv���Uol�4����>7��^�p,�����}�2 ?QH�5a�%�>��#uu�N#�>(��I[��u�aՄ��p�Jo%	�vGc�Z�*��D�k8=2���1�א����/���m��3�v\'�+n�-����+U����:����Sh�|T��	�=k��i������b�N����ܠ����D7_B�{��t�VH����d.� �`5oW#�j"��U�W�7��K��K"�h*A�%<��遆/���XlxV64EB    fa00    16e0n:;��qs����{����Z�u�i�Q�zk@T!>�ZwM	&R	c��%$��T�X�G�⊐K��>!fDuMX�\`Hevud\�!�\�V��V����(��Ԛ<d���[-��(=WZ�g$�I���=sz��I���<b�JY/�]��K����=��?FH�GQ]�M�jr��ow~��RH)	���+��v��-|��W7z �����av��!8@����H��;,Iҍ}X��p�P
c�2�0Da��+ک#�2ƶƨ��n�9O�-�� ��:Uj���e�򜵡�wF�=HZ���� �,�1*���W�e�Z�q�4�'eL�j��Zb�(���q��؜A}Ր���(,;T�'�ǔ�qU-;��){�h����$�Qa���؎|߭��7fסP�q���R)SP>A>O���s4�)�/` �*Ka��`T#U+S�V�5XA�(c����mQ��(��7�n������a���B�[�'</u�|����"����� �z˫1�LV�>]#���l�5P��Qʣ�eIT��L�07��U�>�s��S�h�D�R�ᗡ
��������Cv��I�1����Y�d����p� �%�&Ժp��|�e��u�]i����Ok�������j�ďQ
�ȬeD�#F ��;`R.�d)�!�H�co��aoeX!_`�EzJ��w�ߵ��*x�Ԯ��l�pw��$�,Zz��z���/� ��Yz�����3���X���_\^81���� �Jw��Y��_����Lg�_�&���nJ��'����.�Cv�� $OC���-P	��D����O�׌��C{��1�M���zG����Yn# &q�3$���oԅ���c0���ud/hJ��*�)'��ŚB�c�.��f��1IvhX���A֪v�8�0��^`t(�e��ń�@�jqK$�ٻ�E�O��b�G\[&MH��sd'����+���n��ȳa ��������"3�kX2��s�%�`�RN�;pL#(��Z��p�ݍ�P S�̰�։I.#*κ��D��ƥ���ԗ�@2��l˻w��Cv��uʱ
����Q�ٯ^�H���}�L�3��d�؍�]JpX��]t�vK�ظZI�t�Ծ��j]�����y�j����I�d	BO��Q=W�J��<�hS�x���,�$b�c������k�X����߭:9��3v�Ό&26���7�&
/��7�����9�PFe�ZW�m��6���/�5,}�r>c����uR�ӡ��&r������m�MM��w,ui(|R⫉q�{��F|0ai�
�H�"�����\kٺ\��6����q K'���k�;��P�)�w-|��vdy�]duC�
����{rt�N��2����hO7QҬy��R!��jEhj���u�9&����@V�G���D�"�ĸP}��Ԓ'I����0q�Ö�Sά���7��y@W��H΅?�	�DY��("4fg5Y%߆l�Dz�����1����:��*��z֎�a�x*y�Mn���~dN6d��h]��93�m'��˛����S�
�\G��~f�댿�cƗ�I�h=�R[���W2�!#~t�L�q�ޅ�/@D0l�O�I57�8���qbR6V���Kb�n�C�/l�[�'9(�G�9�c�#1Q��6�8�ɬ����V3 P�l��H�.e���C%g-�ˮ��#�`$������������v���4��kK=q�t
�\��c O����6���W-b:�?�T	5��m[���!W-rD�f����.P���&�T��s��z4�j�,��"B��"�
�F�Ui\��>�����w���1_����&�>�����3��tZt�0f{�[I	#�\C✟&*�7a�����x�'��8���OU$�x��
uJ�zF��Gj3(e�� -�� ��g6�1�S��t�^�\)0�C|��L�Da)\�I��R�ˁ�T~IҰ.�P��l�鳳�6��[�	s��/�n���F]ir��I�eWb�ɬ.v%��5{�����g�
IޣVc�� 7;ڴ�'9�  ݒ�`C��d%mw:��|գ|6>KK�W?
ԟ��x���o��e	���o9nJ5K��`����23�H����1�V�wt��*���ħ���aGc�ӈݾ���!�ɔ�K�$�Jm��~���N�A a�ȷ,u��W(,j���ōXm1��LĚR;�Z1g���;p�H�b�A���i�+-~�)@��7��c��W�{,5l�Hq���׃�-��j���=Bs��dT�V�t}qh�Z4��eY�>-i�����\��0ō�5d˩� x��1 ���~"��0�u�{O/<�8�a����{��UN�v"�B�z#��y�RmĨ��}Y��8�o���w�Ɍ��Ns�[��a��<��麼wo(�2p#��o�Z@O@��6WoU�z���������S��c��N�Ȋ�hrѢ�qfrb|ϴ��1.ru<��<���Uh���0���N�*���znH:�@�G�WH���F���OVTR���.y�$9�	R�(��뽤��M��y]K�g۩4����h%�1�le��ƣ�m�}��Jq�!�=}��8z��Y�X��u��$Bh����F�d6��'KM?�`ЎO%�ʡ=\�@�� /�w�5~�~��C� 
�͠
�aib�{�"`q� m��Rc�����d	�Bd^jz����߱s^w;�>�������&�9�Ź�u�f��� ���m��Az�ꪧ�n�8�ι��N)��3/����A������\�_J&B�߲�|!��%�d5K�k\�A��i�=��5����bÖ�+SK�<#X���j����{��:��F0{���sK�řM}�������i��0��=Z���e�)��ߛ,^�Xa�7�0�NFf@9�Z�!R�ؠ1�"�n=pcY�jIOFz�@��Â!��֘����#h�[�%8���%g���V#��G�O	�U8��[�:��/�!�5N[�&�%{e�`X��6�h�┩FD� �<Eަ"���D;[��E��DB�j�5�Sx���5�BK��,�jw(jc ���g���moj�(���/����������Ip���yI�9�#�V��A�Zs���õ ���C޴��=C��$j����&,�[���B�����(p��]A%5���+ܣ`V��q��E`=f?F��//�d�B�&94���bl��f�(��P �GY�b�4�8xS�ܯ���/�B�+�Ƒ�7�p"k\�hy�e���0L햵�: -�/qD78����Cӻ�+�O4V;���W�\�1��y�Z���ᴽ)��$�Z�0ƹA)���V�UTڴ��.7�rTd� ����ј>_�Hb��E�v�\{ ���5b�0��г�f��C�M����󪖇���|�s
�g"~E���yasB�_s��\/�Ȁ�P���׫sЭ���Ϻ����C��e��JlALIZ�9R}�������#z��e�P6vc�ؖ���5��ڍ1�C3����6C�6+o���]�K�`S�q���R���� �L,(O����Z����󃢈��S�t�#=��:��v �u���QG6)����_�Њ����7�K�aD=#�N� <��A3��附0��$�bnL��dL`Ǭ�m?Rd��i�{IG7������O�GE��SgE���*�oWHg�]!��Op�N$(�a p)\����Y5�y	{2�kC��� P��f\�h�9�P;#�����b�<��ݤ��㜩�ay��Z�Փ�a����F��������w���_���Jt{������\��L��Ɏ�'L��I�W�~��u�#��Ko�V��S�������}˒��7w(f�������"�:�[?M��P�{����g��TL��N"���9�E&:�<������Eʃ<�Dȸ��[������5�wc�纰�i�p\�;��_�Ob���8�P0Jg5H ����@��5��~�;��5y��X��5��q��s��,л�+p�w<E�<biN�#�3��C�.����m��=I�.�Ʉ��� <�75|���UC�8u`.6��";����c*}��##�o_�X�0%��� }}�~�P�: 3�]��Ȅ�p|�S��2�$7a.�A��h,y�����՘�2�T�d�%`C�Rū��5�b�*�[��l�?�~|8��jx}ulx�O��x��G.)���<��Y�+�q�z�0^rr�"F�=��Y��?sB+���ˬ�� oO���x9�G���0g�����>��4$��	#���
����*տَ�6����Mq�&Ə�d[>�0Dz3c��c�����r���{w2Z����tv��5,�&��v�_ �A�%7�9�`{�q��c��ʛú"5��R�0sS$�<��H�1������_ �6���`��L7r�r�,���-Xݞ6�>� ������s�&K��c���R��3Ĭ��
~��ȝ�&;�t��M[>��<S�D���������.%?L!z�r{�u:O�*I);�)�yΊ��D�d9�o�I���8I6@��x���w�Qn�5�=�vWNXL�n��[3FٷhNt����*wd�9t���v���k�R+*^\fz��F�K[p��o�7�ț�+�{*x�%E�QeS�,� D��T�lơ��G t-�m�-�8�&Z-�:U�f��T62�pQ.7��P��A�E�a- ��`}+�NZ|1�it�)���_�����X���i�rOg��z�#m ��e��\����UT�+'TSu]��\������˞Zz#-qr��u�=鲞~ �MI��J�1�C���]��G�t�j���s����w�VE�4�r}����W��������nE�Q��v�[��ʜ{��)R���o��H��Ū�dӝ�2�����*:QnaPb�`�~~�P(��������<F�Wӈ�AC�Z�a"� 1���>C�fx��ڐ��!"P��૳���Ǥ:Z��>c;k�	x�Y��G:k�c3BW��2pf���+�0īahOh�	U����� �p3Sԍ�X�٫��>��XZ�l�s
�������yw����Ӎ��~�ZX�N��r��A.�v���S����{Ӈ��)��פQN����k�Ճ1@�H��H|�X�ߏ�&n.�4����g�"i���co,D���-��c��2"��|Np��?�b?#YK]�e&؏驸�EF@R8`�����A��8h��ʡxd�^��n��tX�2��5K��f���΅��N֥3�ژ(X��V�u�yj<�
{���zqICˇ��Y�Nj��^x}���_1�b:?�7�IeU�+�Wj�cArv鱣s�v�Ng*HbY����CA��F�v���%���~<S��6�(d�>��~R���@|�7_~9�f1j�4�)"�Mc�΋�q�4Q��!~^��������?z�o'�;Q��xp���5�5]�}���x�tM��u7�\��q��H׆�g�IbS~������ �/�(V�T��[L$7uU�l�@�)}F'=_r�f9]>��(M9���A�})`��Ƥ�4��-��_�)�����S����`p���YwUkRɓ���3���+�\�@�H��YVNW�[���?0��qG�E�\gsNxLG}n��L�/��%Ԁ��&
�vA�'X9���Ҏ�8(����ݸjd2���;r����:���_�DXlxV64EB    fa00    1f20� ͭ����0u+���ù�]����+��/����{�yl�[���L��c�f=�-?$�zl������_kȧ�)�ܛ��SGQO��pF	�c���a��6�mo)��鏨��u��<�%���9_�"e�Ѷ�s�[��G�E���MJ�$����͢�T��7���������f��V�(X�D�J��x��:i�E�g�2�3~��������G�I��S�!��y>s�VL��"t[q�(�e�s�8���M5:����+v����{$���|��6���QZ@ӽ�Fϟg��	1�� �^*��:��]��#˹��A�F�i�r������D/��X�B5��=,(��Qg���� #��K[�\i� �gx�>���#l�D!�΀��`��)ԫ_�=�q��Ҷ��e�}��Ϝx�Yd��B�r�cG3��D~jX�.�6X�_N�C�k�ny��"IIR�3_?D	Y���T�)�0M��)�ʮ--���j#H�&#vK�I�;*0�E.���4�����Q�2T�zU��+�_���~�V�3��V�,���*n=`I,zN
�B��Ue�h�bRb��AQ�����5������䊷�X����ɯj��T6H���x��$Ee��T�[wT��̀P��XDl��hE�N���A��έd���A��:G�OQ��DB��3��u�z��|��kJ��K �G�k%�����$7�`:7¿��H�O�ڬ"=��KRՒ�q��/V�n�ox=�24�5v<^^�O�����š-������D1��R����X��hѥFm�܊��)sT�|2��QaLPϩu�o	�W�h僩����JU���}�$����&˶��e�_"��~U=V�(�(�m�
�ަ�Q���#���,�]�SUv��X�3���P{`8[��0����?�%�ő����j�*���S�1f.�$�ˈț]U�?��t9"H�ܬ]��o�>d����<���3�%i
7�XsP��s7@N͉T4��:����L=|,��0����;��L�F����G}p���.x� =$�@ja�e�:�uz��܃�?#��)���pQ���0b����/�x�G�u�{� �|Ʒ��a�O�	��X���a�k5��;CiTɔ��X[����f���uQ$r�e���,jz�/��DS� "
�4F�_У�ք��!��P�Lg��q�-�x�H���jڜR�}�T��G�[z3C@�h�u���u���W�c����ahtb�5
w��
%`��?�j	�Ye�G�:�keH*��j+N�>���6������1��?�U��,vO�dI�6��i
&�o�P��+ YG�m�MB��3�3�2��Y��đo�_�`� �	b,�T����T_��������(������ʌ�V��¸7p�/�W��J|�����h����YB�P�Ҽ�%��(E�U�� ���`��m��Nl����$���u�znr�AP���ݵ��q��n��We�h�Ш�q����s�y�3�^�R�����I��Y�X#9�0���F�f��s���S�4�e"�T��L"��MH�z�NC��b=�Kø���i��oE��������	XS^4i6ʎ6�O�U�@Aq����NB��;��Զ)Sر`�����C��C:}��st����5���-3����7'D��=u����a�f�&T�o�n���ߙ�MC���+Oy�mD�7�2�>DL��M	g��!�9t��M��Q5�*jn�B�m�ˬZ���ϺT HK�A	٘5��0�[82�S_�O[d�]̮.Ǯ����{��ʥ�؋�����P��uwM#�լ���rV���/gVw�������K�]~�iv���c
��c��@�8�RM�\},������ōV�BA�l3r�	�X�$��X�Um�^����ل'����
C*S����n���
= t��H���a�ol���/����VX�>�o���C0���$b�'��ɂ�X7�����]�!5	�}�ż$_��s5��q��Z�#q;�X"�ns�)���v۴I&?MD�c��tal�P��q�O䣎�7(A�,���?�~8�+��v	TK�>,p`��<&��������@�5@A�o��'�<n��y�[�9�?�9�MIU�Z/���F��XO��(hD%"X@����9g�Vy%�������[�"k�tA~��7�%K���gFY'*���U*�Ԃ5�=	 �d?ZB���<�?���6�����ɴc?�ݾ[^/�t"ȁʅ�&��ˢ���iJ����?7E�?[�p�����Vv�%�C/�8�;'h<Fօg��2�u�ĩ��YSΏ�S�X�3,���p�\ѻ�c$B3������EMm�;�v�-Q�����|B��,�:mr^�<W�r��q�P�{3��'�$�H�0ngڼ(����r����hOy��� D|��7��M/���T�aF�E_J��^Ō�:���J��w��4���e�cM�t��Ք�u���I��y>��p��AOU�kG[��`�
nu�D�+wiS>�r��ߣB0GN'Ɩ�´oۺXX^�I[�@v�v�XZ�lɬ�����:WE����9Y���>��]���,�{���9F[���<y�j���ׯ8��w�3�0���z�ơ'j�s`�"7�P�N��H������+����7M�X�p�|>�����(o~
��T;'�h���B@3սU�T��K���b��D��V"'$�:���QrB�X�pʽ�n��w�Ŏ�NM���'}���*;��붫>���Z�Gr�#����p#����Ɉ�zū�C��7z^� %Up�W�	*H
	H\�8�M�E�>���mt@��[�p�L�UՓ�f;`GO��TYx�lK�t�A�"D��9�ж;'�W ���⽏��u�z�߄�f��%�PQ�'����I�c�tES4~<Q�Pޔ�|��{ƣt�M~$�-�<s�mYj�(�.�"�z\'��C�)�a�ݭ�};��Q�F-�p�Jr/h�x��oO����i9���Aʚ�����~���B
�ÐYr܃��(丨!Za�[����Ek�T��o��JO�	J��Q�D�ռ��w�����8���f���eY��f�l�(���I)�e�6�'���cj��#co@�_\v�V�f��"�;|��(��=��ơ��L:?��3� �k�zݝ��ԛ"T�_r���.���0w?=&��N�̏J�n��$-�x�<�����se����'�ԑe5��'�{}�v�(��x0훝���V2*u�q��y���1#?Ĭq�Ӊ�D�1*���'�ra���HڒF.�'�(��)�wD��]Bq\V�tg�!�5���� ����x g�p+B�������n_G�B�i��3o���s�������j�p�1
�~3m�;|�9���s`�#��4�8Win]���PѧJ�&rS-WIB��+�]q̚���?uf00x�,�y=��m�#��(��3���S�+<$�U��ޔ�(�QP<M��C�o��:DH���D&z`�䁅\7�yA��?U8'/�bwq�@�[��(:b�WK�q���U�EX%W]��l��p������UN�e��z�l� ���o�.��o�eQ�J�b��������q ��l���d%������Rn`��R�<X����~QPe��几�&4Z�᱆�����1���5�S�y,��Y�:�T[�>���5����<�Xhd#Sk���}F�n��m��Q�f��&�,�>��{Vx�473|�m������BkN�"&C�M�T�]�sq�!��,��z-՟(3���t#@���/5߅�h�x���/z�R~�F؇jM-&Nkv���7��m`o��W��(�(����k����?>�ϣbS�.�� 8�"�kS@�$��-ydtP�4�2<5����wbeoh.%k��A�aH�L�������%bA�՟�O��+,"�
�+����ȭ|�*BƋ}1��S���:C�P~%��Q�<B�U�'�V͞�\&S��������N׋7�����;���N=N���b��t/���aW�z�����/��)g������N���9�â+ �����K+��ѐ������8��6��&�1���;+#���2��vZ�	���'TH���ћ5(�-�4S�s?	�4i��ӶX���Bi��eX������"�H"@�y�בJ揭,M��sr���u��B����v���ф�w�	=,�#�������)�zU��#���?�����ֺ+X1s�j[���4͇%+��7		P)��[>_aF��T66��`L�ҷ��1	<Iu���F ��'�H���N�Z�~�W/�Z�9/nC�p3[jIއYԳM<ReC���1*D�ķ�h~yf�HU�!��T|�H8L4�i����8y$��_P���R^����:�� ��]���o�#6"z=q��^ay?xk��u(�Y4����d�˺`v�.��\>�RNla[j�T7X�K�+!K������J!-d�CK�g�;K��F[�Κ�z@ 0H�d!`�����*/��������J'�^x�C��E�-HC<���Rp����jH"_���[�1�s�l��5M��'��[�
�Ք�斥��aQY�E���]K�I�o/=+	�|J�#�{ܶ.^QY�'E=w�L������bȺJ���փ��f���t���Ru���+���,����~��0\E
^I׍ŷf�U���t�<�q�ߦ*��j��ǈ0I��o�FE`�7�b�/>��N�B{p)��׵�˨��"#��g����D# ��3E��ǥ$>�b�9�z���fz�V�3d����ŭRN�d��;�H��o=�<B�����sC�4RY�18F	X|�H�Ie���L��>�/�3g�2@�^���7�&�\E8��L8	���MC@���������?7�>��7�,ވ�G<�S%j?�F�ʣe�� �W����6�.
���Yn "@��pǦ�@zȆq��:���ID$��'7�æ�_b"}�W�����e������oɔ*1����~o��G*f{��i�ӣ�[QB�������f5ޖY��m��T�s�z�O-S ��V�`P��C�P�HB�}�OgI4�zk�I�ukRY4����[���Y431;aW?9�� �K/�ry�N/����f���?��m�2@!�sg����i*�|����-p{�eʶ;污v�GN�>ؚ�\$�h�_���7Jb`�/h�����}�2O����:^;'x(��h �V~8�:��{h4&��{_M�O0����Ym6��K���|n���2��+��U���-�E�¨d�CEVtS���	��>���K���,+�GC�h�>��?D�<DN�'4&L����ׅhu5;�i�i�)2���6�+�n��_dJ�L�\o.c@�WTZ�n2�Q�)0�>�5��{J�6[�pҚ��K���AB �������]|�E�9��S�cԽ�d��HC�d�8��[ƛ�����������{b����^��u�Q"�����I/I�۰;��/��a6'�б��>�O�)Ӗ%��;#������x�nMg/f�����k��E��D��jc`��!���}뢄��S�װ&M�Ͼ��Q��T�% 1��ƾ�	����$j/��$,-���U\5uH��$ ��}���v�$O�M������a���J��ſ{+ޑ�՞�ʎ��[V�L�>Ҵ.��DF���������ݩ��MZr��D��=���U������7`�D�ڬ��fzؤ�X�=F�U��䱒uO�x����@2zGYUB>]�=��e�W����KE�e�.'b��z�_UBU�n
��Zr���k7�-���K����	�/��=i��bLAJ����~�)L�3Q0�7��&1�@��96H2�[���u�(�@\ls�\�������f1�Z�2�ƣηH�Gg���nK@̛6���n�a4/:�j�"skA��a�l6�~�:E���z�s��]�,� ��#x?�����f��E+r2SѴ�4j�-��,'N�#wo�:UFx���<��R.�^����0ވ����^p%Q�C�l�ZU����]����\z�(ء� F<�S�p�M�jv��aS1�su؛�G�a���v��9�O���"��Eg��:\�����j��A0�-L�Λ�`���|��`<^�,^�d�#+��*�R�rF1&�l�T���6�ցN2�]2*���{���Nv ��ڐ4A�ۗo:�GBBe���[�-�]5��zo'���.��7%;�����4������PM~0����(�y�Q��+�$��Q�{'W]�ef�\{�xs��p�N������(��|��V�O,��#�E̵�=`���A�q���s�ʻu�R��0��W�s@��b�i���ɯ5�4���U�r!��:����t�[�#�L�j��  �__�����m����VM��H:*�����S��eJ������E�7V<b"�ɨ�1~>`?���2+��qGl����U��B����Qjv��]&��>Y�������N�z��g������n�ߧ��T��� �c�ǅ���w�Qܿ����G�݌�DҶ2��B�qW�k��\?�V����]qA�QQs	�b�|>ݥO������­x}x�ռ���ff~b��ȿ1���'5S�1Wc�͋�K J�(j��^�=uCk����-����FS#C��9R�<�h��n�	���k���kWHP9/�غ��Ixe&�|�q�!NΛ��l�>�r>�aKT�w��m��n��{xL���'�:<
�ڊ)�Q5իz\3i����Y�Co�[W+���p�qc���V��5]V�����N��P�Y�� V�����^Y"-�����6ޏ댱R꺝��T&���_�q)	�����:��t͉ֆv!s����%�sJrx�͕.y��.uR}�����ވx=�˨dG���G"h�"�3S���S�����}�o>j���I> _���\���˥��`�eZc�<+�}y�9']Ev'O�CÔ�\k���Ȯ1���I��K"���cY��ב%|���t���'�sp�I*�Y�ь3dRѢ��K�)iӺ������q.9��+���6d����՟5��MnJJ
.���BK�� I�T.�̢���	�ڈ�[�x���.��?�Tp���Z�O=���RX��{���d�n4#/?���CQ�7i��v;aKw%E<�r���4À�g����"��3o��H�/8�F��p�A�_�C�BwkP�S�p���A��P�`:�����y���VU�b3劣u�AP�g���ۨ2���M���ҭg���n�W>��!k	���a��*�zBem�e�v(5�TO�+3z��T�u:����5k}L=��ߞ�mZxS���RLFs���W�
`1�6
��La�<���	)q@	��
��)P�.yE�h���Xxff�`H�6S�����M��4�rI���;��*��6�ѫ�z��z�4�������Nm�]}+	�D�/�Dg�j-yNe
L�r:�	�ř�
mG���іldu��V8K�s4�9hj���>H�i5
1�叮�{N��H�5���x�����:,힨�E��Y�A�Es��h�vh��#�;�Q�Т����%�������U��SH�>�򚁬ƍ�;G~M	��;�B|��P�D`���g�D	
�U�w�.����}��:rca� 2�WsC@[�K�~WW6�^*̃	���f!jY�D>-�v�]P�C��2OXlxV64EB    a11d    11e01G��ߥ.���Qa�G�Nc��h�2����Ե�)HDC=�уT"4w��DB./��㸀p/����6��6�z��m	������Y�᱀����r!��+�޳a��������{ڝ��ǶV��b�-��uг7����n�K�B�7=����挛��.��>/i9����
��S,�u���06���qd��B﨤�^����OG�,�|�_�Z��{��JҸ%�J	��$�R+��yAP�>ry�)�@`*���a-���-� 9J���4���WFv��𒽶�HQ�����V��6�F��E:�-TWP��Z�m�	�O���a�zo��F���@N�h��gi>��lY��(-�t6H| ��zI�Ĩ�5��lڰ#/o3ˏa��޽�����#2	���E�.��v��L�y�}Qϵ�=�c��t���%�N��l-z��пRV��t� ������%C�~}�{_[�X�^��Ku@ʢ�}?M?���ø6,�~u�xV���W)7�CX\���*�*�o���u�u5c:\�
J1�޳����pR�$�`F��^P2A9���ȃ^=r(⢇�\{���kd�mL��H0��t#0��X���i����C-
��r�z�sٿ�szd��lۥdAJ��(����p�jĕ�n��xP����R� ��[NOA]�Ѻ0�x�Q�Q&�v�ّ/ �"��쁴P����
�qy�B^f��Y���,x����\a���K�[ŝ,
m@��'�
Z���������',:*�Z4Am����v"��Bb_;���zQ�37?��6�G!���8�$.C�咛�S^�Hl�g��s���&N��ދ҈T5�I�~����l�>l����<9�ܼ���LGK�<O������[��]��3����)�O�;�'*R���w	�G"Z�$�/uZ�͙�+�i�����X"k�q�����kG�.�#�&��z��m���cb����Z���kЕ
�,e&Rt��KCsʁ�bp��@HK��u���C�-a��u�"C��V�G-�{\Tͩ ��u+fo���aDGa7ߒ�ǫmf�w��(���	�CRi#�
:7�=-���;Kx��E�|r&�T-��Ϟ@&@<J�r�r1��������F�o
�#T�g�y*q�8fcZ_�/Fz��F
w�6Nz<��������ţ�ߜbc4vX�VMZ�?H=
t4:�h�[�������yfj^��C��cN�@�<�E�J��I�y�2=��V%m91_�G���񅆋6y�~p�����W��v�U�i�����} ��s�|��!q�m=�w�Ё ��A��M�]�N���	�#!��1�����y�0�{bq��׃<�\�l���Nv���A�Y)��o@��!^`��e�[̍3};#���y�[:p����Z!�n�}�{"�m�8{��)c���g\{Ipi�Mw+̌��Ȑ��+t��qPG����<f��A���%�.6��M6g��e��6�No�V�8>-���sf��&�A��Pb5I����,��������u�I��������̅熘D��%I�SS��v�ev�� ������M�7%��R�p@�+��~أz�~�'M�jI�V�v�N�����2\����t�,l������ŉ��}rV��6v�&�ѥ���
;��4-�zы�o]��6���2J�����vP���N���EU�z��k��X2D�3�$T|)�V���T=�jf,�`T�D�~Ҟ����r��h���\�	�V��^����"�1�r�?j�7�5�;՟Ol���ϖ�i�ޖl�ꩠ.�������B)��Q%0�R��������dds���D��� Kg�]����/��+��К�c��oJl��C�꿅J���#�h\F��ɥm�x�<Q��(�"���iX*�m�#����D���)��5�.m�"��t�������c���kOA�v����\�ŃHF��k��o��Q.P��%@1yF�N���~Ed/���z�F؁%G���n��,o7-�L9��g�`m}Ԃ4�nT��|[��o&��ͧ�ė茣$S��}#q�2y�g'���د 2�ib��c�o�)X�I�ZU�5�v�u9�ܜ�t��nE�G�Q�� �U�|��+�y(�|�*z�vQ,(�aV_l,\}hOA|2��֞�-Hj��9�gt�ȁ TI�ĝ�6�������Ć|�����S�/
A��v��]�ڄ�[�����w���9%�Nŀd�#:D#6���G��cQP,TI'Xo��	���k;ք^��Nԗ]/�'<Fg�F���b���	� ��1�1S�nΚ�&���NWk�P�+�t_BQ�^O/��m|q��ස�yj#���BKkw�u�(�$GM�06NB���W���ʪS��6��U"pK�u��/Wa�Y��J۫��i�Eĸ����9���h?#�d-;-4Bų���ZsXX��q�bA�M�i2e,yF����ըR4�EU�����B�ɝ�P��ޕ�Ј$�B��l8�.����r1�VQʐ5���~�T���DL~��JQR��&����R��
�Z�.I��gX����
�.jj�z������9_Ϡ:���n��-�������g������v�H�~�W�s�6��Òx:��Y�.�{I�壾P�U.�����mrna��Pq3�6ͨ�e�������Ж��3����>f��iL�����7�r1	:�p��˂{@�O�'�C
V$�~�pFe,ӂ*GE���;�rg�.4��<�/�ܭmύk�#i�D�Ǫ�Bמf?4@W�<<y�c�R}�����
�2��%f� p7-�i,��q����g�be4�����	K�����(f����I"�L(��h���T.4|�ӄ�pH���#���H]d�Q�IC�u���4.9������3�YH�
o�OB%^�cW�)�.V�T��6��6�
��8
7uP��ؓOs�8���h��>�k�g�	�H?b�;|����y�����Q|�_^�^��=}~8�3�����J?A<�6߮�Ld��G`+p�f]��&>W˨:t������jê_����qR+I9�#�ja�gu�l��FN�9�$ť9`cӇ����ȱ��W��h?���ǙxB�":nZ�9N5��	�i�́f8*f��H��ݬ�.Uz:��]]+G�4����,ё�W�F���X����t݂O�f�w5���iB�༇�?�H�L`c�b�H�5�e�mW�`DOk��p�~�;���DO�S,�
��G�p�Om�uU�\����cX(�g(�U�|�p���~�*g�T���lT��^�a=����%�ME��E;V�RObw�P�����C�SP��ky�>�t����<��/y���'�/��8�TSH_�u�-+@R�TY�Y�������ס#z����[69j.���2 v6������Eb9���UY�t�����X���s0s�$����H���HkT��л���	�.�Hk�����h�'t���c���q�n����u[v �\�#�%ck�b�?���J�r�h���뾰���
�+��SI�U�7�6x��(�\渚��ή��|�f�U���n%P�2m��8�-fف�ۇ�OD��͍;$�N�p���(��*4t��ʷ�5i�c�J���m�z#WӗF�Y�YW�ﲒ+뚢� �Tt��@&%���'T��cty�ä�И������m6Ɋ̙�6��f�Z�_��hd�2��R��˰G���ċEZW�!`fs
1,�y��?�7��$Nz㦯�90����$S}��,Ր���m�2ɜ*f�ir�eX��ӕ��&x$�zŢ����s�IP6K��k8U˿��^��V�n;�.�.��Дt -x0`qw{Z�-W�2����%x6+�	���j�pʎM����UN�>/�����\YA��7�#���α�jJ�쿫WI���C}b��E�W�uF���!\#�8����CWH�� �m�� x:��\Kē� �$���,��z�dX�C��F��Sr�&y�<�`�*@�;'�ϜA1����+?<�����yvC��R�,�{��>�����9lN0��Ccl�F��LF�R�6S*zȱL�UI0�����-n���_�U���{�[�a ����OquC^�D��Th�y�r�dnzfW����ݬ�$m�z�?!j��1]'D�}�U��J$y�F�u!Κӑ]�y�ɑ
�Pi]̈́�:JfP?�ص�>�'�'� ߔ8�:z7�� �c���К8i���\ɋ��rD�E�E��/vS�E`�j�JW�Uo��T�<�d�R�Խt�,���!��p�q6T���^{�6}��wm���ؐ�W�0�3����]d~����$�"{��k��oM1�_ok�����_��Pto]3,�
Z��t2)�6Y*��6@�zݓ��*���OD�ޞ��/%�qv���VWhv�#`���c