XlxV64EB    39cd     f10:U���H�ش�!$�������?����+�#|��Cc���#���-�b�i��ϻl�z��D ~�|K��thɀ}*�L���f��y��<��;�`�����h�؏?�H�����*����P��,��n{��/�B�Y�ê'<}�9W5f��0�{5��S�7-4���Ys�:2��w�J�������e�8�Q#��]3P_��'�c�(d͛�@��  l%��zc+�g���@�3O�w+
���|H$�`q$7���<���+w������? �aoN*����x��)V�NN��r�K���!UvGj���n�R�c�b0��R���\ڊ#�����F�j���Dp(V��_Z��(o��AdZAn�eZ.5�_$�K��+�y��rL=��ƣ��c�X��Z<�ʸ|���xu�d���Þ����m���A�&����}�M�1P]�>�_3o�Ŵ�F�d�C���>��+��pZ��#S��ƞ�mQ��tF�ұ�����d8pr��l!�_~t��rj��\���8�7�A�x1�Y�'lT�_���K�T񼭭�Fe�Y�H���qx��4�@
�z8i���0�v<�i�`9��g�)}��H ����5e,ܨ���q7=�N=�g��k��d�;�4�F&�	T�B23�~�%�!�,���N.	���߃�	Æړ��Pk(V�&���g��	{x3딤�!BC��/������2c7�QYl�(����iT�&4�~��7d/a-hZ�i��M����ӱ"�~�:��ױ��b(&M��^o�@$�����&#�	i�"�d�;���e��E@�/<�z$rT�
8E��{��n.����h+���h�$��==(��K��z:8&��P�����8U�ɂ��%�!���"E�y}��Zo'���]ՇY��M#�cc���
��K]6 셈F\�7�BL(ܢ���S+���J�(�ZL�L�!��9��~�f�{��KR����赒���@"�/�O��?��"b#|;�\rLR	�m\��L�I�ۥ�%�)�u�"��v���1L�f�h\��8�`�r
�#Dz��ާ��/����Bd�'Pd��_+�X�� V�ŧ�z�=dY��Z�sJ՗��+�f%:��2��G��v�R�u��N1o/��Z�����Ζ�N�e��7s�V{�����^wWB��=� �-�Ȟ����Ty�ڢ�S��8�Q<�=�t��kx�ޓ��{^�x�b���/d����?f�]��OdǶX���$9[J�S���`�%>T�;��J�vJ��{`�]0J;�k���c�u<0ܽTL�	�Nb�����<��R�g`�L-U�Oę�96 �I��oL��ގ�T��wC
��?�R�b�?W�g�ae/����w.qo�/��a�O 2x�e�݌�K�`�>ΡE)����0=�uH�����ў)�=.lR�a����^B��-��'��sCTtx�� �}�\ƘϬ��=��v���HD)*Cy�p��!J!:��<�0W����F8tw$XcBAU��\��#�u=�_�C���Y櫫��)n8Me���$���u>:��y,�!L�W8�T�Z ҂��
��P��t�D��AWq�S+a��I��m��Z �>fה�t��!��`&���1s�	�L�/ߦ=�n�#G����6�����#�{�����F#�~@�RFS�L7[L�4T,����s���Q�uO�ߧ��r|��@���C�{�O����f�@� Q���>�.���[���(��$���F���m�j{�ڕ�7<�����ے�;�ya<T����~��4_�L�} t1F}����*`��g��l1�S=�7#j����1�.�5_~�
�u�"�λ���_� �����H#/�:A;�*�a���<����KW{���-��H�6����x�b��8���#,�N"��P`�ξR�QԽ7�5�}n��\?��MoI��,�*|��fb����|l�7>v����?v����J�ڋ���7���Q���ɸ�O�}-u��-x>������P���;�k��<�����������>j�a�%u����=Zmހ�lc�P�ub��v�Kx��.\�k6�a���NSq�c�UD�B���mE��3qf`M���n�#&����L8R�ņ�G���0B4��Cֺ��7�b_�ILc����o�H�VEޓD@=�ǃ	z�9�ʠ©E^�=JX̶�Jl�_&o�Eju@���*�߁Þ\�B�����6E(�;��IFTW���)�[,F�s��/���;�X����������t5W���`a��|3*���^e͐l��|�aR���~�w�v㭣í���}��P����Yv�v�E���!|����Mn�iJZZ���Bt�/h���k#M�}��G�Ih^�T�	zF�YGD�]���g:���wb�Ñ�ߖْ����K�M='����0�K
��P	邃-0#��"�X�_0��uy�(��B7�7Dq$9tmj��`V8S_�����0qE�A��4(�a:�T�d�Fn��ԭs�c�2%�:��2�d��g�����9� XU�}M��z^�.gr����Kr��D�������N�Q���@�:U���?.�����m�'�ky���#!ɥ-����i��0��&_GF�8K;q�j����Xq��X�X�����4=U��tO�V-zVf �����K���@��ƤN�Z��u|��r,��ɤ�k/��T��ժ�^�_��B�y�G��ug7��k�gH��qc;��S�`��@q����|JB*Ф�J8)Q)���"	�k҆����t���;:7��!,�}fw�7�?��=��T�P1F����?�/�����E�욊W+5gq<�B��|�@z:��b{@��g��la:�Ւ<T�]��J��ål�y%g��:��6^��z]!�*w�,Ț윂"O5�:��@���t��u[���Z�W��6�����hy&��uT-����=k<�a�Ã���w�j܅��="8wkXX(V��$�Il���z��f6t:X��_v��S�	�.���5� �����lΈ�=���쀖ٽ�����I�����e]4�`��D�x!p��]	���T��moB�r���V�g��r#6q5��.�4sj(ʨ���G�����t�/��IXD;�?��Z%,��78�J�yg��!�_�l�[\�qX 7b�Q^�����!ɹѡdP�#�l�╉�&�8hՉb���^��~{���2����yr�\=>�m@ݗӤt���!�:�f�D++#c]֑��ZK��N�@�ɤ��>���e�q+FZ��B�#ت��gsN�E|�C\��=H���=|�@|0����П�4���t�{z�!�2 ��pJ�^c�g���g�j���Q��!�0���pU�#���l�&	jh,��l%��D�X�kT��Љ(�����q��M��Y������m�@�띗\���Cm��7e-�vG�������	Ch��,W��(�=� �ksl������T>>��3z�{��cn�ˣ
��>��pZj�J��^��W����B&U�o�z��:�ɔ��W���h��T4��\�>M��]�&*��
	�����&�oI���֩J7`�� %|�N��t��k�ؖ1-�*(�l?���OyO�?8�{P<5|A�S��P]��_
,����k��%?�Ȓl0<K�O�e�E,���L�y?(i�w��� 'UG���FA�1~��p$���d%S�ƴ����