XlxV64EB    2706     b70�.U)Qp�iD4pVCu��r��F���V��G_��Y�������O8/�;T�Y79_L��]e�����lx�;�r��A��<'ѵ�� �INz�ѿ�Y��9�54s����)e0�Đd�hv3��Ɲ^V&���T��8<���Z�1z��^�Fb�)�@�2���'d��4�SA�C4i�Љ�%��d��c$��^A�eX���\�F��A���.4��L]�s�5�����7ɻҎ�$<��:�k	|Tǡ	7���VQ-\d��E��t��j$�\ԣ/�d�%��˖!>�}�3?N��|����]��
#Y���fF�#$֠
9��t����h�Z{�>���)k�&qr)���Okِ"\+a՟�W�xHk�NDR��x�H	��Ox��������PbIR���C��J�2��U��h�P0�_�(Dƣ�1ae��S�V��S�c<>3�a7))�k�d�͜��<�u@�L�o�y�V��,[�-㴀 ?�U�2�(����'X���(��D���ں[Xs��֟^$� ��Q��"?X��7��� �%����%R��QHc�szY%	�\�_��hܰU�X!��aݢ�+�5���6�I�?Hb\\��5�Ը:%~UT�����`]���O*��#
�G~0���ϐi��"�@%�!��Q��&i��ύgr����/��<�L�bǞD��BH-q�K8���Y���	ΜAg�NY��+�{�FVj�7���.�> $�U9�����v���<\�u��͟�L�{zm��N���4�;���T/�x�k@uQW�eZx7����t�J�{=�oH���խ�Z�Y �����T�ӛP80��)�1�a�j�'~Ə1�J9�����b>|��F������b5�A� �4�jF����8	�Ƚn��5q�H@@�'�5�݁�p�b���o��,�as�&Ӭ8D��K��լ��/��ٍ�b>܋�I�~�ֆ�=�rS*%��6�-3�|W=нC���/��x?��戆���܃d��{U6���T�����'�bȌKm���ʣ�V���^�'x�Q���OAqB��`].C+���JJ�,)��.�Z^O6�\A[���"`�K,{��C	����
�i�2�i��İ��/��0�ڙ�˾�����S�K~������a�Z�+��r<
-��; ��X��Hv��Gj,�i96*e����1j\,qܺB���}�G�������~vE҄��q�8�밴9�3y9�����T�����bo�M���҃���f���5ix�YDBh`��,y~�Wѕ_30���(�B����Jݏ�W@g����޶�\6Y͌$Y�|�H��[U�4���>"���%��\�GB�C�xj&9��Q�		�gR����|r�����:9�4��iZ	���+҇w-�A��T�n�}Nכ|��:�1h�
L�h�a0��������	��"�-����-];�9'�sCL�z>���Y��(7��\zv����H����<�M���^�D���4� ��Nܡ.�3
�]�'�/�2��鹧�v�6_`Q^��jhd�>�嵘0������x(=
Tq�]g��=�&��J����oq����{�.����1C��g�t!���!�68]�p�\��O��r�X�n�y����P��|���i�/c$�ǝied@�3�Z�	U ��l4���t���(ۼ"l��U�)A�J1�2�W9A��J���{q�� �F'��-�,~��q^̉ 6���T�z*v�uX���^q%����=&��Ř`��]�x��)�<d��'���?RBp� yq����Co0F�܄��x�^5�yG�pQ�tw�(��Wȭpp_.�Ԫ��a�$�sFkOHā5�%O~'4��/.`����挖��m�'5Ϫ A��6&{��eH��Z��s"n��E��jf�-�?��LS������l�}�����X	�H�az'C6g ��~�d���"����n��3n��� \0Eb���*1����J��׽aY����k7u�=5c��)��T�2���dN�m�*���3��<�_��,a_u?ݞ$��	$
cc)�3�4��xHs�%��iƜ[$茢��羗C��x�%,�JޚrښU���g����tqLvs��Lo�$�v��|h�����T������&�
������tƚ�Ֆb�R���S}�֙�`'R�����b�[[<�R��N.d�/UT3��W9 \T^.e9]�����
���!9�ps!
���}V��peq�4X��L����'��:
<!���j�	?@7w\�C��YfeaV�ѝ9�t��� zEe�~`�pa�K�7 bG�%_�sG��S��G�p������#V;���]����we9�9z���>J�v�d�y3�F3�OlX�����.{p�[����O�R���K|II�Qy��i��1.�����Z�=%t�=��p�'8�%L�9p�
�z�c�ŭ��\*ֹW�0�&,/���_�B'����uP��<ϝ��82� \�X�b�1��Vb�:l�غ&�u8���ZEU��Q�	e�@����lHR�h\0��������[r���f�g��\�۽�#t�	�q�V��j�=���0���t�RR�,��+��~!y/��9�4uİ����^�����>��C��t�s�j�76�x!U򬖖'RW���;�U��#���U�%r�ra���%�V\ڹ��%Wƶ�~Z���<���#H��kjAVH��!�Vq�3O��DE�r���z
������4w��"��3�KO��[�g��1C�� �"��e�&�pI�Z	��U*X��|�	�[rc��δV�/A�O}bm�L�x�>�a��l��g5Ǐto��F$��z��