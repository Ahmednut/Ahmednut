XlxV64EB    5716    1300��� ���n�g}�:΂�����1xq耬��%�4T+��#́q�A�6J��kX����Zu�H˾�S�"5"��"�F���]��EφDI���6�������&��7e���{��#R�R�IPO�{�A-��o���j��s����%	KW��H4
ǀ��)Vw��l"Nɛ��qCJSJ��(�ɒ�����&�#n>��T��_w���H9�0��p��"�zf������9B�(���=�E��K �5Kd���9���)��Q|Io�ջ+H��xkV����3k�LY[��x-��W!�Zf�tVxj����|�'��h]˷���O��ȳ�|�`��gZ;*�H`��N��Wg2�|�Ƚ�M�'�{�	J� ��is_��S�[(�A�[�Z�Fdӹ����TքC�3)F=lr�aHl\��|��I�O3�L����ƽٌ�aR̕�*-��ɇ>eV�����E���b�`I;�
)�}"HAev��ݍ�E/^��[̈���O�B�`W"SѪ�jU�\X����͟��s��U�6�>f� G��������T�.6t=+�14h�%���A��U�232=-��ռ��y0���L[V=�"���N��g[��w�Oþ�T�X*U��=�^�eA��Ԯ�8��V�>�h���$�T3���@����N��:$�O�a%jP5���r}2 �@h9@��9��>��|k���W����F)��*c�1�?	!M�٢��6X��-Yd*y����_ѓꐰ�5$���(ݐ&�����=+��A�$��o�7��ӭ|����EJD*%a;��0J�>�<T�EJ;n�r�)��|�"���)��N��-�yy��+`�ܙ@�{�qrL�D���p�S���U������;;I�g��������uC6�B�Gս[���n��G������CJ����ۗ5n큹���Q�\_���B{KōC>q��^q{����(7�p��i�:���:��o8*(w��9L|����E9�Z�R��+fP-�DB"��*��H|D���� ?iU.$�Jz�~������ƳA�-����]�A��[/5ko�Cr���X?d��R)A_�9h��U�)�u�i�,	�bg�ݚ��7h��qo���o�<�A^�N��g�`�s#��Ǘfo6�4�1�ƨ<��Q����){���� ~�
�0\��-W��l�.Zdk���/���ul֓@��a�E���B��h����.�RR��@|R�(ȟ�����x����9Ի���Ì��D��3a�i�;�8 6����:u���2�h���%�C����p:B�W�7��d���ĩX��ěta��M������9�܇@���w�L���s�N�66��.P��<�U�Wf���d�e�#���q!0+Vh��
/;R�`�KU�kʋ���O|ѿ/�Lؙ�g� �[��^r�2ap�:��*��2����&�4V14�������
C!.��#�c!���玒q�7���֩i�>��؞H�B������x�e̝�"�*Q1��'��E3��ο��Z:B���|T�;nP~7�{��8� ��Aֲ^--pt1�0�	fA�+�:w�0۹���(��i (���n��i��T��a�Km�o�'��Y&Sy$��~��gsr,+�����B?���!��"5��)#�bz�H���{�a2L�U����N�ĝ�m�}�_�N�K�g�;�ĨW�h�M�!p EN�2b�ǈ�m���G*j�c��HV�z k >��F�!�q�K���>;l���
����r�}a�x�͹waw�Y�:η�;��ǁ�za>r�BW%+3ȸ���ĲI}=�K	�ƱF0�F*ޑ��\h	>/���*�6ܮ�ٞ���C�[��kn�'S�Y�'T̓g�Y7b;Q�M��-q���T�q�F�!�k�wh�:z�C?��R
����¾|[��1h��%�Y`��ƿle�8��o�nE/[��S6u1��fݍ�N?3�X�g�~�>���di`�C^[�#^gP#�%baaO���9�Qlq-2����0ʯz��B'�m����*
�'K^ {�Pp�Gd�W�X�d"�����1�K�K��5����yּU@u$AD��9oMCޑ������!R�g�7q?��sU�X�%�} .7�����q��&�YU=y����Nnc��ɻ��,I(���	��@�s�Lsw*�T��tᢛ�{�۳��Kw�®���*�B}W!q ��{���,Rx�}����q; <��4HN����Tuؓ�b�.�4,�y�*�KJ�]�V��
_���n�2���NJ�Ιj���:S���"�BH��?��;(�}�dn�Sh��Y�8�l�Ą��ώ�5]�Х��2��18T�)0�T���]���il716���'�5��O�'I(�{| �Y<��9��F�ƪ������\�fG_�}�Wޗ*WJ��"n�4�o�
2hS�8݂O����B�4v^����^j|���/�V�	���¡�4�Z�����=C�W��@S��f�<����p�Yo��~�\j������ ^�(�>٩�g�$���J�A\-�0v���m�6�i�B�_�9DK��Q/p�pR��R�Q���j�Q�%�Y�k�\�a�>&�eQu:�!B綢��lsg���p�ģ%��g��g��dS���9`� �ڪ�HOA�d믕��Q�!6_ė��pkZ=��@ZD���.?YP*�պTj]P�i��t��X�2 � �r�}�a8gĔ�����-�M��� �G���D~�����t#rG`_B�g�4�]�3��MW�Y��_�@�7���0I�/Mo�G+��X����>tq#�(�D4����n�ڻ�׹X)
�kc���0xu_ٛ����]��=�����<�H��������le���#_�TP�-;�:�M���j�W��1d=��j~`����s9U�r��xf�i5ˬ(�����"?�NR<������D��6%��wi�������
�ϛ��_��ZKU`�'S �ҷ�6
E�/YA��j(�n7~6\�Ehe̂D�DӚF���%b�ub�����J���< �+�V��C2ȑ8�KjR��,��s��(�f��Il�̏1�s	�> X�-Nˁ��l������f���2Y�3�B�*�a6�����~��*�3��؃��Y쑵F�|XnjL�s���>�m�<���ul�	��7#cn�%x� J���i�0�!����_���7"�W��Gr�J���s4y�U�<����m�z5��8#Ko���]x��-�10-7��iK�ɰ�?\�m�r���TB@9�l_��*W�x�(�K�,�`-2j����L��Cg��M%яyͼ��'��������T�>�M'�S���e��с��Y&:�t����ŋVT}��n
���.�:��Sy˄5�мn �@�,�Ë����j`
���D�~��$v�Sb(�+��'��8���r_�5ZT������(=�f��+��������n�H�m���<F��n�zR����Q����+S�-�j�&2�ȻE~+,'9��Kq7ƾ���i�ٴ��Qm\7��敏�+S�K�-�f����SQ�R}��0�@t�#��:��'ًf�v�޺�^���tZL���7~����;��)F��iػ���o�>�X(	RQ&�@vW��X���Y8�Gm&��?�<o-���R'd�).��Z��6V$��a(�Dj�����a���Nν͸UU�[A{�3����Q�՗����T�=�ȃ��lS3Lz���&������RPnx�`�$��}'�cU�e�lfj_z(�	*�|PZ�u ��\��RI�G瘐��l+��Xn�r�c2!�H^�D!Ag�l�W��+�r�g��Jr��aR�˃##��W�Q��0�p�ņ���1��n�y\��簳�l��S�\)�c����=Sa3�U���D(�j������HUGMP���M�F������
�c�%��z��B��[�ʪ�Ee���p"8r<O���&~Z��9�tZ|�+� #�U@>Qq[g1��[k�[�D�!�*��ۋc���^�fj�>/��yq��o]'����`�KуP�}��,�#F�w{��o?W�_�J|�7���v�2�Ԧ��G�kܭ7�T. 	)���q�F�:������{��$٠%J��}��n�;��O�%�!�ZR��U���'r.>����͡�rr�zܵ�W�$�y���n9GK��;�i����C{k5_4��u��G=�7"²O����vYh��wG�~ϣ��˂��,��c�m8]�����SB��mJ&���9�$�|�`h��$��T�F�7m�u�xl����w��y�����ȝ�� G��7
@��% ���Y��a*TWd0�1�S��[�� �ћ�G�U�Q����7�� ����F��Q�9u��{r��˝
SQ���T��%���96����(X-S�0�}�t��$��F�h9s�5�x�`ʛ�]�C�NJ��*�2._���,�9�˼�vG�9dm�e����d4r�PT�]2�Ś�9�h� ����#J%��~W�|bQ�ĸp~��2,���h����a!�O�����~�ܨ�S8��2��f�8�3!ֻ�����Q��m�e���溒��"�,���|V���:M��4#Jڜ,���K|��u���bBfj�Z�Պ�S@��!���{an�l-D,�B������<	cf�7&tƳ�ڎf����v�ef�\ ��)���Te���` t�}��pR~y�VDT����Rz��ӂs�%�(-���Al�C