XlxV64EB    2279     b00HcxF �]\5Bm)O�WZ�i~���@f �{�쏧e ���>1uO�P5�s�bMۼ���Ԗ�C��f`
$��3��迠��$��ί@C��0����N�o�g�q�5�hr���f������1�,���������<��*�c�v7���5���ryl@��6$9]�Mz1�&	m��^}7FH�t�7����#�h+�,�V��[�X�0i��ø��\&m�B�Pjۢ`�V���$��#��b�b4�`n�U�3N)ł�+b^x�p�++��e,�x��.��Jw����z�����
��ӂ��w�d0S�?Ժ��ӌ�4�iS���`�E��;Ď��da�2!������E
���mq��϶.�bE�M�G����*&^�0�?#�9��'��+�jPI��!�(v�@�VS�N2.+���!��0>��������Z�OhЎ�]�-kx�:�U@�������j7|�[��q��Q���]c����5;�	��舴�����6�M�mi�{��.uK/r$�5 +���|�D�#l�s��6}N4�,%�H�v�;��9�^aྗ`�?V� S��3RT��
��P��d����m~ei�WZ�=ӳ��ߎ\���ʹ~wP5x�S��r5�a��V4�y��A��`)ǓLJ|�e��[�\q�]Ԕ�J �u��2Na��f��08���0�u�_����O�jy?���^��A}���i$�
Y�c�#�����{s�#8䲘4dAFo��������Kmw*����g��^&�9��BO����ı�'�����B����>���u���C+@*�u��}0s:?�����W��� 9��'�})Jś^��Ĕ��*A�7��<�M[�͡���$��B\��J�y�f �1+`��VU�B�[��c#�\��R�ީ8�4'x�`�=b?�(%ɚ�yΏu��w�>gA�Gé�7Ń��ۚ��t3+7�㗐�,�5u0«���MQ��ЕI^��憛��j��M%��I*l��fR]���~�*�(�r�7:��֩>�^��oϪC�p�;��p݃S�ç��f�_2�BE���S��_ǽ����v���o���w���E��EkY@��>d��"�Ĉ��1mA���R��pU�2���=��\�SZ� -*߅ֹ|�!y�ج�������b���/�) �˷�D	+���P�6�^7�+��؄�Pc�%Ԫ��~�24�@B�_G� �#��{�7�ר&h8�H(�.���	��t=LlV�;� �f���̖��l$�lWi���n�#ģ܁J��f:͘�XO=P��'p{
&ᤘ�Ǉ�}P��Jy]�,d��8�&���')x�$[��x����fR�T�Ƌ��}�<����zӎ�5v'2~�@+��]�K��@s�H�Ie�p�"����r]SP�|G�dS�q�E�y���}�Z��nv��6�`Fc.�M�ͪ��_i��)݃v(c?��`�+"Z�6��T� e�x3]��]��J���A�"�0wM�I�̈́;��b#_wL6���Ӵ�b�Q4�!���s2��1e�A�Rm#���܅����m���6��9�S�d�֮���Ooy�k��;;��N<�|.T�*��E0-K���"�g����j޴'h�l|#�f����ڤl�@�����rQ�諆AC�r}3~�;B]wjg_�/�A�`�2εlb�/�����5�
�O�D1�z=<�s��*��7�C�?��rt�
��������v���2��3N����M��cg	�d�X�� �^�Y{i��)���ḫ��c�=O�C�CM�7@�폳@2o�⵼{R(���a��Y�!io����--�sm��i\�p'�J|�/ضi�����E���N���(sn7�(�;-�����v�A_{gЧU
�G�k"L吊��Ю�?0��Z����k����$�݋�d	��<!���X�E��B��:V�����[�^y���h��$=q��Dx�O8���Z�^��ZA�C7fP+�Ĕ����,��j.�`�e����F+&��)���Pjx�5�N.��{���?po*���3BJ^�CPmd0�YG+����r7��U@	��z�n�Һu�]��b=*��f��kV��~�}Pj�N*������{-0P��>��c%D����ܭ߻�Q��`��wrp����$�x(��n~�#��Znr�4��*w��|��w*iP�T^g�n4?k�H���q���H,�d�Em�-p�n�K�M�OF���,r�0MF\)����̈��W,���1�9q�!�ꊙ�-�Rcs����>S�[�ͨ���R�{a�/qO� ���r�H�r�r?ɽ`���̬�|�3+�͹�'8"^�#e.u�=1����!�VW#�t���
l~��
����>��T���Q��� C/Y�h>Z-��e�7�(X`p�d���F�xC���ƶ��Ϝ1�۔S��)O�L�[�$3@�>�M1�[�`� y���B(�5���O����p��/D:.�J�G�B9�>�qY��r��_�v���d	|�Hș�V]�THT�稞��%�b����Ir�$��T����/r�ǂ$DKv,2i,
 FG�9X	���� :���}B�	�ʭRď�����gF$���ޘ~_�.x�?�]]��ú�Q#�?�}׽���?B�hh7�AIky��{� m(C�(i��)q9ނ���Pq*�P�_���N����$�zZ�AN�8&�d�jƃw%�!�%<"*��@�F�8