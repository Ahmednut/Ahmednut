XlxV64EB    fa00    2f00$�<��a�_�f�c�Q�zL��ߊS���>r����m��R�l�}���4�;���߽4�f������sh��Ħ��6P���=��5�V��l�ҭ�r:��vo���&y���@��"�^��w'U0�Wc"���;2���܏P�O/�%چ7��嫗�P����;�E�$2�svB�� �'C�m3��~7g��A���A��Ԃ��LL��#���k,��G�~i�B�5����&�Hu��6Ղ���帢�YU�4{�Y�;�ˢ����+�5[n����/����~!��l�!P{R�_�� B{���;���.�j���f�����Y�z�q���Hȝ�/�JG#�_Q^�z��kSٺ��Y/u�ߝޢw���V��,]و��i���'w��q���v�R�%�y
��o�*f�"�$�h�̟��X4�zG��G[�zd��P|C|���q\�z&�c������j���.oH����?��e�R$4�b��\��wra'���s�J�a:xk�Q��5<
��	x��W�����/���5���w>�J�]{�D�;.�,����K�a	T1=.�}�*>L�w;{\�(��F�5XŹL�1�0�ܑ��J.�doUe��S�����ȮhB`��)g!C5�H�:�-?|�M�)�����^���!3n맪���M/�Î��-rJyْ-q5������j�R�o&�����(����3��'H��+�U�h����0P ��wXe)3"��?����	+�Yhc�;��6li��T	-�Wo{6�l�&J�eb����p�XbL������h��q���S/~m֭j��=
��.�sf��G�C����N7�-��f��p�Frz�t�"�v�'(	��zm~�6�;_����'8>�7נuC+e�g���*���r	JŢ���=f�K}C�~:?�I:D����ݪV����d
q���������?���2�DW��\hq�z�������Ba5Aio5�~WA�"o>	�@������&Ri*�j�<�k;=�a�o�;7Ј�j�QF瑕��se�����o���7��������_ +u����G��(�|E��܎	F#!E�#M���a6��Ǽ��l�0��7���X��c�3�n�,�r�=�*��}^�����Kз>L�`i����9�q�dgJmǿ���9��a�� �s��J�G�R��Y�qN�_&��E�_O����O�f�����`����N�\p���5Ѿn��uà�yA�'��U�tz����C�is^؈����%� hq���-���l8s�&�P�䑮��aSf�D}��$��_��|ɓ]�^4ǎ�\�EZ���aIA�2�8>y*�|�ڽ�{o�tI��G��q#aL�V��F�#B��M���z�!o�vtF��k�H�[�-'Ց�ЃN.�_��Q玒_M���?8�`�1�@����U��&����|x�=>/��Z |b5t4B����0���@?��CT}����v���^��̌)���t@X�����S��$�=�'_Smf�'K�����C���qY��ÏO���>�}^��li�Zj��iQ�`Gi�mCX�Ձ.Qn�Xx���bE7�9�N�;E����1���m�̬e�YeLO)�`X^��l�Z�Z
�=W)����,�q�ķ;�7UJ�=E�ӌz&774'��AL�����hs��i<m�U�7F��*�~u*o���o:l9Õ�~�n{�n_�[�M�w�_y��� ��!��K���m������c訙��4><�%�����)o��-._�#��k������>�}�Mp3G�o���g6��!���Jj����$3�O≆���sXA��.4~�/A���\�vq�6�[(�7�e�v�ؐ~;��r���P�6�D�+a͞g�@�L�P�*B�"g�mt	u�U�R�*���R�]��#(l�֒�%�zA�E������t����|һ�A��V����Ԟ�ʀ�x�Q9�3��=s��,�9�����Hćז�+�e�.`�&�!�f��i-�Ӕ�w�o����ԛ�!�B�#\���/.���F�s����q��x8��9�MFE�L�7�jè�;���&G����F�$�5v\э*�(�<��4Q�;�<8&�o%aJ
��R�ڲ\������J&b�q�A��,��#.eKk�A��V���`�x
,/�Iԅ�	g�Ǝ�e����U���c�������va��6���֋���Oa���V�����I�q3��Z�(R5[VP�V���`j`8P-���.4�Xb���%9W�Wʧ���]��t�l�M^~�R'�M�4*g=��)���UC��JS��ԣ6m٬�g��qb��4k�K�V�:��}e��@�=p��.s���JVg�	�Y�v�W-N|V�V��w�z�Q�2M���~��	��ciC��e��4^�W8��5��o�����5@qF.�؋O̖2��C�Y��	y����qq?�f�tP�u
�ho�p3`�����M;�f�L+F����>��7c�
�P'���Zja�������'��t�wuht�y
0������4�v�бyަ�Q��\E>�h2٠�n���Ȝz���e�#�(vt���fD�[��U��1]=SWt����4������-l$պ�c����.�Yqf��Ɲ��Zz餙|z'�,��ˤ'�/߷�v>�']���f9/����rv{���A�Ƨ[S|��$p�>>l��>�0b�nN0 �$�<�����d���y�7#�A�����+���A�i�$����_�w~�����Ӊ���\�0�����T謌����2����ӌ��!���Ia�����wGzo��s�e��i0P'S�V|1o�u\��jO�s,\j���>D�����~�Ʊ��U݋ {�Wje��\�&�7�
�=	���w��ٴ���h���&2����u��I�x���}^vѽX:
T����̥0{t͚C`��b�~d��֨������n@IUi�����ߨ���#�idM�Io�楰|HǨ�Z�є�۶�.as��I���^Y�����ڂ*�<	m+�6���C��e��#�q��d�#
F��^����������)ը�L��R���Ժ�=d��k�C��	0�H��_DNPX]�
3�@n�>��O���W>w�f�R�I�=/�Ǚ~YA�zt�[�L߬����k����p�� )P��l�i4�'&�m~%s��V�q �����|P�~J����7Ig +wW��7�$��ڃ���6�P̔+*$��|[v����0�{�"�.k�� ���P�QV\(3���(�K>kZ��~�e�a���BA�;;���8�}S	.����(���F5���۽B�\�j�l��'�ݑX�|\���2����_ݿI����E����X4wC�)k�"-�O��赸�B~�:\�ov�(���#J�ˈ���*tUdR $�����������Ex��~���~VI�{_%�k���e;�c��Hw����Œ��������T�m��J����kB�����(�c{��篃���'�ǧ�N�`丌e6Ͽ�2{4L�4�{�SXQ���N�v�ܮ=6ڽQXY�?��1�7�O)����n����LM7�m�Z�y��`k��1�De�ةK�&��3o/b�M
D0!0U~��)��:#�8D3��ZBlD5@e�%�n��5�ի>����;=Ǭ�|q�a�\�Q;��u�M�?��;R������KO�<��vhW�4���gt�2��R'�"Wi	Ю�7�����]F�ř���M`Ě)����W �^z�m\��y���D��P�
qԗR�̵^�8:�v8��Z���/��Ai^m@J3��P������R1BK�s#����#�T~�ash|�z��.��ix�`&S�o����;V��c\iO�����p4τC�Hc����c��4�1lʍ��"00�U;�W�u1���m��ld�d��:i����D/௠�t����S@��\M+�	��U�L���au�䟡�-�E����T4/D�B�8�]1�z@���GVϖ���=R�����:T�ѽٖ�$��.�� *ܗ;�t1�H"; |� �v������v��vn*xG��T�����XG#:��K��[�8�7Z��]I��U�7]�;��.E�Mlt�1�aÒ�7�'�Ϟ�Ή��`�ɠ3��'���1���Zi��=��M��@L�՚I?t�V�]�P�m�?��2�fiT�������j�|��K�<j���S��\S�������������������9kT?��栗r6Yh������T�a]=5d��$Շ)��ӣ�2����b�S�j���wJ&տF�8.��B���i�����I�J�(
�
��5�e��\~�}�f���vG�w�"ˁ��άb���"8�)F�k��.�l��#�F�������J�,� ��d���IWƴ�Z�������R|������`���ӭ�M9Z�V���\�H�U�\���*J�υ�L.(���ْ�D:��8 �V�H�􉦹�RR�s�?KK�9�P����5G
T����tR98�n��mh��ϲ�12>|��S^��J����"�I7V�-�m�ء�����Q�� �TV����\�P�@���Aj7o �̳�&�Fo5ۈ��A��Lқa�޾|eu��1
�L94�)��/L��m$3�D�zn_.���'J�t�?�'�
��u?-#X�P��2f Zi��*x���2���\rO^Qvz��E���Zs`ح��ɭ)����;���B������1�0	��u*՜'�� �Ce�hui�r%��Կ=���{����B���b�g@���Q�^�/:�U`����=��NWɟ�i^��>N����\�{�q/�/?;�i�7>l쏈�x�J����~�(c7��&&��6ZZlo�#�}�X5R���J�k�M�?r�S�A�@UE���wY�VvZ�&�y����4�c��䋽���)���GuH��q�!�W��]W����J�E�Jr�>�V���/��\��'�X�?���$�;2x,'JH�*�Z{F��7�G�8�oT�J��#�\O7"��9R'�ц�#֜�� ��o"$R�W0O�f��m� o��1'��h��3Q��kҘ�"�amαS,��s(��&PmcL�WRe�ł�a>�O_"R�g�p��%	�`� �eN��Y�b�)Q�� (��2N
�2uJvrLÀc/YG����[\zM�1.X�oi�d�guw��+0���Hz��%bWQ���su�i�g�/U�0����M�|O���2߷��j���ACYkk�.w`�*ۼQ��X�0��ޜ�82��O^�M/Xc��6_�0�U}p��k��W������0�8�B�����׿��A	��w�� ��!���B�IvMz����7V�PO6�L�����a�Ѻ���.`'����t#I_`8�Z�m�ұ͵ѧs J�J�o����e�<D4�S)ڱ������Q�η�ǻ�����q��/�g�0G��f��&��.���a�Z�����[������jr<�+,�Ļ���\�BM�9S휽��4ZZ��0�����8��tk��圉d�;�F��Q!�l�:&g�P��)� �7���a=�bZ�hv�6����;3蝿����o[�˖�w�KU�_͍mp.m8�:V���l. ��~_��y�8��2a�އ���_m��NN
��f�R9��}!���5�Z��'_�_�d�u`�ٕO��LXT�V�Ȝj������Bi=aw9�7�#8�	x(���]Ɔz������._
�hXV�%���L5�=v�.ޓ%��Y��Y�	�f�l�Ԩ K��#tS@�冀�֒�,�)c���eE;�~ӀT8��#ZE�wr��eSS힧*Q��I�ܨ�|�(����D$���G։�m�V'G�z��H��s�~Cb)�ĕ��垫#,.{�i��vA'��0f��W��B�n���A�p�G���0��8���f�S�&,��9���H�Q�*&ʏ��*�����mw���&0�!nŁ��Az��C ����_�=QVu��~	v�-�x/j#�rI}O�*3�B�?u���P'q��ީ��\nW�Ƿ��D�&�.����> �!n�����Z���R�Bc��F��eG�kߑ�b�(y-�R$z"��[٥pv� %i<Z��ͨ���B�(aL�~=M�;Y���s��gI��iOǌ����x��{�Х�<�6�7�GQ1�ɲ�;��)��������k��ԞRM�R���I�ɇ@��rY����,6H~�Z����r��G�M�Fw[惋��/G'�0Fh~{0/+l��LM���jhTz�Pձ�e�+������70�✧�mA��G%im�5g����ƫ	|�&կ/j���r���b��*�s8D��2^�ͼ�נ�b����Hc�>�}V�R~�HX���:r���2� a�E*� ���&�@8VYN��4V�9���G�d����3z�¨3��G����v���G5�%(�@����Y��l��`�s;�f�:���ٯ���=�Uh-g�3��-�'�&(�C�#�}0畚��flG��~�L�Uvt����K��L��\qvxC�b�w:R���N�Ik���Q�2\U�N�Sx@N��y������sF��
�D�0/|N��%�t���kv4�����N����ʯC���ܞ��mD��ʨGeU)��d3���*��wcm�Ąp�����l$Tvs�u�s�Q�,J�� $�*Px�� ٠F��Π�!�FD�1��ε�E���2�t[T�����GBl�|��$�r�A��*��.�]%&J�cc!ɍB���I�mBQJ�3�5��)ü���_Xv���_��ax���O�ّ���F�O�A��9~���o�=t��.✜���<�"@c+w1��F���N��E x[� ���A�
���(�*\��㍾��[U�gl�P�$,oAA�ۙ'���ʠ��8�i���)ZNGU�oBp67~܅����<s�K�䜟p��T|u���$�B�|�d�b ���۫k�!�."�9ɰ�j�~Q���tF�%H�h42���ONT�x�4.���ŭ5�6�R����|��}�!c�X����0\]��������70�NJ{9��؜��,K��8����-�:����Ew���]}�,5�6��(y��;y��s��3ȵ�YG��<v	 sx�/YY<X;x�i��b"��/<X�B�x�%w����Q�\��qa�.�~dے��6n�2����>�q�t���':�Z*] ���q���r��<���I��(��n��m>�~]��Fev�L2)�[5r,�}��04��N�yh�r��6� yEOK�%��}��f��q�W�=�\w�[ṋQ�h����2�I<@b~�F��EV\0%̸j�VN�(Nmy5�o�n�p�
@s��)�#B�UPລ�����o��p������0���?YI����wW��O��<�z��X)[g��'Ak(���8gI��L5��Ech�i�U���2E��|��9�o�&�;��dv��t�~�T+1	��'�}�LÂ3c,������sldgd��a�ϟ5�X�6ۭ����P����U�;�[��aس����\�o9}mA5�n�Y��|�ޓ�	���%j��,��Ǧj%��$ʓ�i�)~JY����<-$D�F80X��50�Rw5��;��L�����'A܃g**5okl�a��ޓ��O���l$026��3-����\�cp�}�	�\��DG��ݍ���}��̺�6	�V�^(!�O�LL]�lՌSh����z���ﷴ>��;)���!�87.�Wy3��d^p��'Y�	��ą�(��Ajn"��K�b�S�>��m��>Z����\N�|z�@X2�F�\�-��g�;���u?��W�MU�A��7��{�T����x\����t�1f/.^U���b��Kp4��2�wl�$�8ԅ�'�P,6�)�c	��Y>��?r^�{���(q�gC�����~�����9�B�b���gA�޻'����Dە�۴+�<����Uf�7�:۪��oڻqy�YSŴqIT�w�BA�
�0���3����&L�C�;>6��B�.���2�7p�~ p0�p[!x@t~f�ki��b;�%�XG ߸I���Pf�ߨ"�Uz�J��~�)�cu��*Yɸ�OQ�� &�L�X!�6�l�0�g���H�O�62y�Y%[W��!�|.����95h�����1���,Պ@���5!%j��Ź,��. n�Z��z]�}dI��paÜ��_YM�z3k>�|Eu����b�H�6݉���.�!+�c�ky�>���!����2�QT7J���-ǵ	�g`Pʥ$�eR������+DPͳ<�~�lV(s2U���hWr�������==U|��UhhǊ󸜏�
��E�(H�	��� V�ɦs�g2UH��n�LS�bַ��m&f#��38}�� �zu>��P��zd���U�����{�H'���Rkg���ݙ\�RE<���q�5�R��7��_�rE�jÀ������ڣ.�		i��Y��n; 1Z#�R���� �pm�"2t������5ke4�w��D�!q�o~�=c��ఖE��y���j�kb~}��g�H7s6��k�%�b�ڹnEd*R$��4�X�7w�X��,�?t�qS�WN�NMpg"+߳pɨxTO/?��w����]�e~�ϟ�x�Pu���T7��c���ҟD5�4��B�����n�W^mU����pH�2��j��A�ƌʎ�}��
5�
����X&�㊈�'���V�9��[~�� ���ș�[�/r��́��= J�Zy�	[��Dl����K�3^��աɰ>b��P�&��u�S�|��U���6�RW��8o����vb"� �r�
H���en���#���px{�Rw!k�Ƽ�i�{�I��a���.[e���Sh�1
wu�L�|���eC��J�!a,aw���V����@�L@�Wg���&�+� ��T��0�|�ɷ�~�_��	��L����В�����6?\�12Wּ� ���3�g�ZW�Q��:3�����3��f�0�ݟ�[�,$"']V�v�t����W��ʐ2p�K1ﯶ0V�⇱�T07w�F������Qh�C�&{b�)��]n�ߣ�p���=�O�BYȁ�R�h4V9���aACJ־�o��g�w8�Q!�X
�dpH+�.٦Y�&v��"se_@��*u�� \��>=�E& ���4@�)7��V1�	�)�[>J�!z�^�1I��I6{Ty��k� ҈{;}^� ��|����Fd�ЈWt�P2 �1�Q�˽4�X�r8�X����ّ�,�P�LyL��$�M5q���0�K<��io/v4��/:��`)��)�#q���������l���G�؊&�oZ$i��ʯ�W�ք�&�۰�Ct��Pq0H߰j�
���f� N��E�����2Ft��Ѓ?ۃVA�����>��N�s�I�֞�%�D$l��Bcq�l���K�m�u�Ï��;B^!�X�l!y�_�CT��}dݵ�@�:��1��ܲ�>�Ç�ۮ��XM ��2�9�|帜�ԛ���� �eH��z8����-%���E�9�d ��L+�����_i6Q�_�_B�tW���9�@$�!Ԁg���h(�Oo$F@c# �����rN[&�=�B2#љ���V8X��Tw���/H��F��Ly�
�]���GX.GVa�7O��F���z��f�c
B_�pԄ�bMR4��gB��i�^T�Ċ9�U
����a�ŵ��c�71Ec
:? W� �t��2r��T[4Z#f�/5m��k��<ԅ��{0Oߊ���@�{�M�j�`�']ӓ&�;�L�Ȧ�
-ChNHx�x�$|�1���ԣ+�/��[t�)"F#g�x�����5*�|u��R����:�|�g�z5�h���{�ni#�9�Y�y6�8km��^�_a�c�6�a��~�f��x�Y�a���_ E�4�\�E�	�<\H ڍ������C�i:
�%����o�"͌:c������F�d&�Y���/�Gܳ�tV.F�a�u�G>�k�� � �5'�bnb���
�m�om-�'{{��=zCF=!�����.;㇀��������:�m��V���+n�0�f��,$Z�Cg����o<?�߄ڱ�U�ȱ��x�ft�Ќ�Pj���L�R��t���V?��No�=
v�N�IH��<�����5�՟�'g��+�	�-��Ht�9˵	��귴���(Z4�����	��M�(!� �!�i<�������ư���N7�ewjSX!?S�bK�'S�=�H�߄n`����c7�Ƶ�F�����`,�Ff�ͧMth�!N�)�9�#�gVD!�]�|H�N�%KR	CP���Pې�!���:$g&�e���뇫�j��=�yR�.��VZ�B'.X.bmY����3'}�Y�;w<ď���I����l�O��O�`ڨ/��u������4��?�Yl�7���LV����7g�n �S�ޙ{Y���	�<T-JL��at��_����?|2����,��CI|�R�BB�}�����rԻ�ۃR;�P�t�r��%�f~��]{���;��(���p�|�,�4Qy����O���������m��n&�7hf�:#���k�?CXGq�1T�d��<
��-�<M����|�̓�������/3/�Z�h�f돵�º�*�<�bН�pƘ����I@�\N��4�gr�Md�ﴓ���%�������#xP��0tw�Y��#��뚐�.��]@g�1���h�bԅR�x�.G׫�zGL�(o�A��s�:ZbvZ�.�gܪ��⑥�$DxI��#��g��<�T���d�<ƾ($��Ҳ^r�P��`B�At���Ӏb3�*�z�G�Q��,t ��&��9Jf�ë��_qi���x��²JZ�wժ��m�j�c�btGҁ�eƓx�XH�t��Ӏ�E�>���˧��?�ψ^��v�γS�j��w���e�N�R6t��E��7x��Pe��n�0\im]H� �^�~g�ݾM!I@�jn(��|�BZ��΃A�~���\�Z-�ގt��WE<��+�Q��0o��΍6\*��G���	
��h8�yn�W����!zBR#R��/L�HB�".l#� kf�s�h��H�m���ޙ�9���}|� �Nʛ�8�������'�*�r�Q��zd�E�%��������IF��6{�J�@K���v$�Z�=���.�^�d�Z�z&j}���N�H���KD�`��jÅ��Z�Q��/�%a��̽�:�I%�?�"Y8�~���Z�cHY1؏|�2�\S�:�}u�h������V�en! p:ƉA;6��՝'��y���%��'���o�Le
�N1f$�A��q&61tN,.KV���ku��F<Q�U�m��/�:p$��]R�$��P��hR&��Xu�s'�Lf��j3���!��l�}veO�7�pQ��k�R�7�ZT0c6�K���A�4!�Ϳj���pKT�Dv��7Ao_��<{JU��x�ٿh�X&|n|��U&j�|'xbW�
mF�q}$��ԡ���v|X�R�#��A����Jg:״1�$�sl����I}�u���XlxV64EB    c30d    1fd0�_E]դ%t�+G�Q2R��}_�LH�']����"mSN2\���\��sj ����J(o��*�89��a�T'�`��c�$b"%��� �X�`]�QK?U��`	��!�,�t�]%\Q�go���ǿ����ak�qA�Ç���[_I�������=N�lE�+����:��[��1�>�_����ML��}��a+��g,�Q�!N�rf"vi�!lc*�m'`߉�$̼Mi����f $fK�F�U.t�bX��#�R���TY���L]@*��<��x���#R�C�����CջCZNG9�2��}��v���-�� ��~Q����N	�(L{9�}��װkϘǳC@��C��
�� 粵$�%i@i�%��~>�K?�R�+���A�f?�|�G��A��&is��s��c�\9��Y`�¡ߴ�������}垫Gl�W�t�p��e��o��,�EO�>��Tg	&;�,�Y/��J��� z~��%� �i��&�����$q�����=?'�9�[u�����ʧ&�7�^Г6���_>���O���kmKw���P�Ț)x2����fX٪D�J���n��՚I�4Q�E�d�-4����A����L�߫hu���z�خi�xŇml�@������X���C��h��3%�S#���w�<������C�pbo}'߈Q9��yH�L��B� �kg��ZHΛ!EVYL��글��E�wK�����erq*���L��\�n!S��[���~8s�y�*r��jx�����O������-���"3���"d���ը�3�������1:Ucmz����;@����=[�VJb�MFW�0<T��Ĝ!Ú�b��S�k3r�ǆ�@� _Dwډ%5ɨ���Ja*ĜC9V���26y;�ǛJ-yd�y�9ɡ��:����_)�s�E��r���l2�qSfH;i/��z�$Q��6BA��a�v���L\��uU$&�4ߏ���Q�D4�'v|褺bE>�^
�>��8��=�`2�v	�J�; �ꐼW�uҩ��lG����4�\�[�\�ں�~gc>�;�̞���{�$�����&��0Y��QIaCo�,$�M�0��t�>_�Y�����L7�bNn��LV���k�#�Zx��J�\�й��ͳv}�QmV���] �JXH��Y��9Y~i�2�I����V b�tv��A��㭀7{����������h\|�]e�=Eߟ��a)�+O��[msȏ��9�3E��3�=2O~;-�S�6j�|4�vR�\Q�&\��NPDG�����Ø���Uom�ޅ��� Z�E�OD6��2LP�m)�������<0�1������
=�\�a?Ƃ�K\��`�1���~���ZW��*%w9̀�&�2o���x��Շ�kg�kR(8ʲ�#nV�r@冟39���s�ئ��A��V�\ۅ+˳�X��Q!�.@��d23�Oz�*��CQ�`>��jl�0,���'�ך(��ɏ�+�	��}��^(:++��(�83I&́�����@|R�����6
�C7'���L��\�C�h��ڳ�V�$X��f,%|Zx��3��iݩ⠻�I�N~��9�wO%B�A�@xVj�F��,�e��u�>yN��M�Q���=6�ۖvͲtO�EVf�;��i���!�-���ܥ�A1S��Hm(��B��Z:�d�Z~TaBݽ!!�ِ���1�
T����_}	h6���L���H�%a	�ń�,SDωz,��ȵ�H��ڕ'巅-���I������W��@V�'3k���NEIL�w�mż�M�"K�F>�S�	�z�הJ�-ЧT�ݗ��i�8��r3Wu��7�7.����gmg������p�͍>"��Ъe��;�T ,Il?m�*z�����&c�˘��p|�ڼ���G��'��|.���u���1�	��p G&���
M#<������e��$�tF���z��eux�S*��/��6�F0'�å�T� V��P��c��v��r��F�I�eoS�C�7'��Ϩ��L}<B� Q�Q3E�\�m�`Sm�{)ȹ@������=�q��]0�Q�a���cie/Ƕ:o����[H=18n��W�$0F+�֞"!���A��%��+��O E��]Y���iGӇp��
�+���u���,�Z���L�%ta��r�IZ1.�jB�T�4+gDj�=�N���D�@���X4^*9�yr���G�������p�hu�-3g�&N^P���w��63�I�_?*!�R� }ǐ8Ǡr�,�G;氮?��:wFg}Bl|��L/���;�����J�)��̘>�)�*��'G����1�	<Wԃ��좣��H����F"�iK��t�#K�����x?�r(�jn���z�Zd�W����B�N�`���} ���ֶZal��'{�&J7���'��g+I=S��돎�&� �jٷ�,R�x��l�Hf�O��?L��%Ϻ���#n�ʱ��P��Q�V\� .I/���)Ϣ΅��(��i�M	�����8ف����X�8��B���*LC<Wz<�qT���S�2!�ܶ��qej�"��4��.�Y&��i��8�-�F�O}j�HY�n��*�_��6�V�8��
��g���g�8P2�-O���-s�Tm�娍�m�ul�Ñ���J�Md�m�Nc�87/���L�>e�Z�Ӑn�n����K�(�,G��OglM�Nڸ��'ڵyЦ�����r¢U,#�G��>c�d�\���u�`ZϠX����-�ዶ����q��V&��c��k�m�k��YW��Nl?��e�<ȄS������C>Ӵ�y�7�hh��S�b���0? DUS��Ӈuj���3�@��Cj �#�(u�EN"J��n�ڷQ�~Pkb���fk�%��/�4���d-�E,`H���X�����S�6(@i�k���rk�?�ѨV�!����B���.� =�J�`�@.�Iķ�k;�{Wtm`#ܞ	F�m}�$[�(ԍ�%��\�	43S [�s��'a�
���(�kD�E/������&1lg���I*o��NQ2�ְ���ƚG��asw4)�7/���O��T�2&7�o&h�5�5e�)/���h����R�Jz6���N!���U���#��OW�0���e�" ,]�C����弎���ͺ%jC>JQ̭�.&H��Ѩ��+�GuJ2w�iiט�ms�Hؖy,6���ȕ�v&�J�ڶ=
�L�@�C�N�m�3�_`#u���ק_��\��92��?���%ܿ�a+�����r�㦩G��hQ���x�<�o9_۱�#�ja(7�j#�S��jj]і�0PA�v_�A+���o�n��\�\RVC�at�����-����]K���t��0=�j���h#�zj�b�� �#%Jz:v⼿�tq|$P�́΢o�NBJ�ȓ��4��1"0���ă3/w��F Yv�<�ȶ����C���<*v�G��zŪ6�GF9y���u�z�ܼ�P���Z��"pI��)+�$��u8I�xA�2s������"O�=j��LÝĲ��*�y�-"���&h>+��.�&��Ի�4ؽ�y5�9$����j)�Ϟ��X Ǭ,vN�	�*�����fN;X�6'?{½R�۞T�0�F��i��D��� �U�2���^�rW'\�&��N�C�1y���\V�Ȫ�G�N�S���".jϰF�p
5բ�t�
�2��W=�F'Tlc��B���K_��}����O��@��\��ta��0�v���e�����u�@���sx,g7�y���4���Q�ak(?�.E��"��;�7AX�� �;��Oq������T�t�������f<�����wiJ�y|���ŊH�hXm�O�f���&���'w�7MC[���/�j�V���_�Ĥ�������L�I�����,:k�݂]�����+} ��c�e���}_	\�+J;P��DB��1��W�����|��Lj�.X��A��(q%��r�v	��������X�Z؄m]�Q�!�b��s[����T�A�>Z7:��=�݅�J���/�S>�����JȪ��?���.���ul��皽��@���]`����z��Pk�8�xg�����_����x��uT���[�8�#��QZ�t�'OI�����*�O��B�U������MG�Qg�#Tj�[��`�Hz����-SV{B��*���Ťu�}\v�@r�I{I�X�'*�]�΋C��bi�W�C�2й�{��p&�R�W3�Y��Ԙ���7ʹ�Mh$qwQ*Orrl1��	q��z���Μ�+�å���(�s�MՆ7�~� �_���^W)�����c�XB���[��Mm;��s��"�}��{��*7p��9�*�ө��#��}�®�L�<$"��l��tq�Q�����$��$4��r����1��J�Qlg �#9���Uٌ7��~7ٴ�T0��v��[���=ޚ����p0�Qb3ϔ�
�N}Y���_7$տq��� �\�����g�a��Wl�>��I�Nqa�=�cO�W��:'��b��dk�sKt�������<֭�?<fp�QrJ��u��h���Vj*#Z�%{<)�(Ԅy�K����i�u�u���bw֌2�j���	��x���C��F����*��H�ܺ�ɷ�zb�a�y��;���8ZQ�����<�K�o�u�r�,X�Z�1�0�,o�/w`$ޯ�B��d�s��K��e?2?hl� 7F�4BE���>.7�|�[*?������?��_W�S����h�E�v$]�Y���V�"-�5���y��Z��l���$:2)�hܣ2Ч{-�T9�!�IG�#��H0�[ނT%	A9��p��#�;�J^�Y)�H{aWqoF4`ˮ���Ǚf�7A�aEe'�ڵ����I���MȷsakJ�����VI��Z����$����GP?3�Ѐ�R����s�)GQ��耛�h���>P�a���0J?b�&.��i��R��+�8�Q���S)���y�_��Gt;�-��/�"u"�/���a��@�wT<�y�Ȟ�a>|�lz��@��T~��_J���q�'��F��?���S����p�9��e`��vf��Q^�pk �e�%�S��k|�DK�4�4��8}��Ie���a ��ƸlDc�ϓ껪�5���3u��d�7���g�.���#(�?<~03���a�e2ǋ�.��R�199��|vW7��v�o�;$^���1�yH��.:�.)^tM��{~W3;��s���� ֹ}yI%��^ո��P"A��Z�bbLkJ�Ųf�;�˼HSz88]����E��,��)� �ģ[0f�,�>���j
62�(�֌Q�������/�U�ɢ�����]�kBw7��e�Ƌ�uf	\6�~�����x���+/4m~z����ś=����y���#\�G<o��r~O�&���;��G҄a�om�SX'��E� \pk�2B	��lA�.��h��\L��	�A������)u������#-"�z:,8���z�.�������AO5z̃ǵ��A/PP���r�����K֛�cK���T�Q�W����\&�Y!�^v̺�Agğ��������z8���M ���3Y��O���@�����h0Z�h�zr����0�S{hC@W�{;{����L��M� �+[�o����wYꞨVc��`y)E�1���q�OF�.���5x�_��������Ф�-�+ V�r���.�#�STt��(���[���?�uM�0�Au���2�಩��A�3wA��D��+.G�Ld�=�=�S���3�c�Wv=����@�Ͳ�6��׍�<�D�E�B��VÏ� �9(V=�\����H;;�����aHq6�U�N0�H��#��U��v��Ɔj�3]<���=K3F�;�����]�Ё�m�����*�'�\�Vb��9����,������?�R��_I��i�Y9��X�8���N؝�E��:O�)���{:����hMe���EZ�^z�z��	cb�m	q��� y�'ؑ�[1a�b�[�ߵ���Gz��/�`�����Ѯ5���B\>ʰ���87�;_��|d�������ù����a�H����@�@WBi`fS���2�/N�n�#]�F�2\��s���N<�� !�����������w�*߶�0r _�q$:[706w�JK�h�VBY� ��i`�e L����9w�� i�M�5Ǯ85���6弧�Aף��y���d�:Vbn�p�ޔ�F�������Uvɾ@�qGPI�zf�x�(���b��0�W�}m ����7�Q�b���b�P��Y7���]uU^�͛��R�5� ����ҭ���&�w|r��V|�̅P=�r1��hv�yǼ���J<'����
�{�ӝ1M�H�(\ʠ6�CA�i�9g�.Z.Lu<��ς*S����H�GI��mĊ�Bv+pNn<��}3}]��-g�b�J�Й<��A�7!IV��ͧ.�U�����W|�N}�az�$�c�iFߩVX�����B�k��J��Ƨc���d�[|-�#B-�jrB0��6�/�/=<������\L��#��Y�ؕ��-tGˆT,ز�4+��4�~=�z�B�F)�6z����{����|�%�����)eń��ҵ|�T]fޢ�xTw.��W�#D�O��\���)��z���ܒ�Dڋ��;6A&^��%�e}{"�̆�m6��z3�O�=�c}��$���Z��l�0��˕��P-�l�3E+F�m�?�Q��nY8и�]��-���Z`��o�T�M�JHe'2^3�A�!<��ڲ�F��� 1m����T��<�w"����"S�:��a�W0����z�jf
}Y���>�@����j)6���/�mgb~pRƝ���Ǚd�1E���/ v��{�E��v1��w�7SD����)yG$�?=/b�/$���1�����(���V�Lwp�j��k<���������.Њ�-?��{�\A������z�_���W��roJ	�}���j��A�x0���[x��gu��:�EW�kc[�҄m�_-��8����H�N�+�%�+k:�
��9�������U8Pf�Pme�։�X�`���G��v&:������PD�2��>yW?­
��&8����J�_^��'\;c�7�M�N�6MrpP�����k�ԅ�G��o^0�z$D�/�@� �j�W�q�ޅ�JQΫ�uNS��P��ٱ^
��ո�#�ehy56bg��ؚ���Xm�3�a��h���g�s֑%C����O�#������'���LVd"����2���G�"��S��u]zi�Z"�[#��X+�R�첒�#T��)�	�51�衟kٹ���@���&���z�.����j�<ؽP�{��� ,��?�2�5���R+G@����9�ց�.FU8�v������dt/>��HK�Q���jQ�]����&���/d$�
��$�m9!|td��$���i�2Ί��(����^�=N�N_b���=Яa_�~A�\�A��ÖF�HcJ�0:�NY�ÒC_��a&�%�#k�����}��JD4�����v����1g�*�,N�y��$EތC

����
�8��ߴe+��������e��E�؆�m����Sk��a�Ow ��xT��(k���+jc.Y�	�5�5��gSQ�)��N��%�D�����5a�����A0\'�ĭ���Q}p�g. ��]��'�I$�(�9X�F�\J@<k4-m��a3o�	��^�X+ʖґCP��Y� ���N�}�u
º��C�Wy�-��	<�S�Eb�����ō ���%yQ�|$�ӊ��V�O	���A�Jݪz��3��X��P�2ք�B�w~rY�����9�C71q����)�AƁ���{SP�����(*���I���a5ak_���~Ԝ��(V`��2�