XlxV64EB    3466     e50������l�rd�L��f�XaTɂ���io=���7`K䙷�,�>*��|��sZ$��0yjUm)着�x��3�ui/A�a%�K�=m�3��X:lʧ�[p�m�_��gA�[�f/�60�d���q�l���【w�}U���h�ka�~q��Ғ��>�	�����yޯE�!��5�*)+�S�t2wk5�G3��ҡ���7]��RY �(o�ذ�5���mw���"��|�y�(uLo�ڡc�kn�3DĎT����
ߨJ\ō�%+�
�Y{�;�����t�# ��$̛�ֳ��Dl˵�-S�&y��Zl�2(F\2`����8��D����	`9�zw�9������K��$k�<"�-�G����;�un=�8�l��������_��X#�sV�5��pn[����@���^@� �{XZ0��p�S!�5F$���:����� �� ��F�� �A�쁾�ov[v)��Cv�-"2���� OL�v\Ei��!����g�ݖ�|�_�m�; 1�5w�Yn�*1�,Y[�m�')~
s�RbeCtai�G��[��u�޻��z! �{M�$I����"�C|�Z��4�>���g8����0KY�x�ૃU5�&�s������}|�� Um�$�C�,u[�g� �Y�,G�A������U�W�Ѱ0���՞��@~6
aX��-/���J t��w���uk���ppQ�Yv�������g�@�4���ZU�2%xm ��'y��2]ʯ⦦`,'�T�Y�`T����?��Ҍ��jQ>����C��J���c�
��I�@�щg�~z��)�E-Lx�)���cW�P@;=g"��QW��c�ŷL�Ĭ�����9���@��Z�6;�Y&D���������s�u���y}{�����R�������q_f^���]J��|��c�ouq!�ݠ�6�P�ze�][J����ӟ,��TA�
��@m\v'�xG�P�e��Qկ�f�W����pnZ�]�pƷ��߅J�ަ�8��M&�C�vx�6B"ȳ�����}��=I\����ϳ��S�tiP����O���Yi��j-�&��sǗ)�?{��:<�^j��Ҭ~M��K>B��y(��H0��:�z��q�Y�00��Tj5I@2׎/+�~ƴe��l[�3
����}U����4.�NLb ޜ�{ı�ˁ��B��#�!)������nǹZ~(���a*{��"����NΟ�j�i�И����GX{�삱��3�6;��c�۳A��v�f��Y'y&X¿B�<o�W�a
MBSg]�%z�����n�v;�2�'`�w�;�<�_	��פ㔅�����]5ԝ�O|�Ğ�n*��>8}�-�x/�\({��h��� Ӥv���	�"�D���+�O6�k�7�d	}�%��~�R���������pӫ���L�q&_�!���+G�;2.��.��wpԫ�޶��q��7y��]u��!�@/�[2O�m��U��B�&
���Q���T��Ⳁ����<�e��n��:y�x�J���F*O1x�՛<�>iT��[#/,vIPx,���� �M4�}ث�V�Ų��D������r�*��J���[V�0��fd��	k�wo�� {DV�H0�qwh�9�*L�CB׺�.�f-�H�O[��%��^�î��C���Q�	��5KI(@�m��T�ط�/��DBX4��%��5)W��v<(�N��T�~C��޿�HL�X Бg�~��R���a3��ب�j�d�u�Y�Su���{b���aY�5����B�X<�F
QwN�;��dG����yV����pH-R�z�Jt�=����Q5l�ӥ|��V�����V�M�@�b�U���54?Y��iSޜ�5�S���;&d����7hs](qZS�����k�#`N�'��$����F��Q6��P�3��Bc���<9�F壜a3AJ8U0S���`��I�/n� ����"z�L��3�ΧƯ��5+P��m�J�s��Aȥz�F�k���lB1Qi`���E���7���6��1E�fu>E��G�A/���];�j����K'��G�ݴ4��j�^�ϔ���1��~Qlծ����r����!�R�[G�\U���u�!r9C�g�x���z>�	.rn���5o��{��R0$�A�O�5H�>�� 7�H
����R�1 =����x��J�6�4LAD������V_�ҌӔ3~�.�2��l��D*���P S{Z\̣�2�?�#ѨWV٥C�Ì��w�5�8��Z��7h��[
�M{d\��μgy�0�^`�f��� Os�1�/J�w-�Ñz��u,�u��1�.v�/o<#����y��j{	}lc�bP��GH�u�ڗR�#��O��'��[n���~I��Ʋ�c�Q��12�6K���#���9�X)T�*^�-/�J'O�R�A�L�gz�d1^'���FM�U�j�ζ"��,B�ڽ��p��:b>��-ϴ�o�uUnh?�
$�{��殏��:sq_�����x%��ٴ���L|��X)���\���u��ۋ�3���6���s c��E�q��:��*O
e��R��;�����v����w�>Q�?�|�< ���68-ٓN<�*����P������K28�܇SP�眏\�CA�C�� "���l��ĩ��%-!lkW��z �~K��������x�C�Wy��<��0S�N=��h��o�6[�O=�����=�_jF�{���!�h�R)�V[�8�"@��Q-�S�����#N���wm�K>��{�Ҋ)¬!�4�$��E+h���`����ȁ�ï�t�g�ʜ��*�������	yb�\@jؘpV#xWb��6������N�w�P�CA#��`�cqEۘ�A��w(��*�x��}�Zj��w��+�?���ײ�,���'���0ʿ�/�����;�R�Wv�G�M5��@�P�����R��xbᷲ0�.$���:��x�du�탁���j�%F��i�gqv-�-�W��~;w=��a�XS�!!EPz&l+���]=�<G��g���P���AN=�DJ����"�=��=�;�T%�}�C� C'Ɣ\6���9�yL�OF�:�X�B2'����n�Q��p+��'���<6a�2b�p�!�/Y���X� a���b�"���~����,4�4��eY���VK�1�qF#�
KKA���y٪���r�B>-�^P��8�����w2E<�V���gܰg�'Y'���:�y$U����
��+�f��,��|���Z�}���B��x��U�vw�:$�鵻�T;�� ����ҍ�&�l`j�9}6�l��kc|Yzz�ǿM^�ޒ���J[�5�ݨ����}�?#�࠮gP^�h��n�W=��3`I �Xm���Dl8�+��~�2��#O)���qw
U9|�:Z��э�4����!����˹��34_�O�슜�-��Ω�5Z�g�P�)��,j���K��V��#s&�7�������^ІH�&�H�Du�S�ep"%�!����YN�3�ĭ@��'[H�B�Z�3�cZ