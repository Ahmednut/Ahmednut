XlxV64EB    2118     a70�+�qɗ�5��}���?� }���G왝I�m�@��๜&!V��q�Y���7��wZn�H��W߫�T�H�P�d�>����o��)Z���	�AgɃ�n����G�*HGz�ȭEX���$5Y�<��EՅ)�6^����4H1�d1���\N���9h^7���%�/
�dN��3hR-yC�pA'g%y)���jd�-��/���{����]9Dw�X�(G-��]���A��QS���$u-K�I�L:���z�%���`b
�ƴFZ��`(����|t��"u�?:�.X��H�Ԃ���[����J&X��7_���.��B�y����+��7�R�D�0���Cnd�H��Pτ�YE�t����z�^��rQ��:A0"�
�l6�?&���ZαnW[���k�%��q<�6�-_�k4���&���q�p���j��e$��.��x���8A4�(��%��-:ᓹ.x�(^���&z2���/V�ͱK���9�z'���1Ҝ�}�6�u�2����%��=�%�Y+�k�\�&j���{[���<7샺�)4�1����0�8b����t�#���?����`��Ƥ\��ti�jjfw�D*w�|�$�`n�Ж2���I.�}f9э�d��D(�i�v+�?���O��ЧP�6f����i��������D>���j�'?.���ٮ:������g~ɑ�va�`SFH�GH�Y�~�P�Ml��p\@���񘣦�C��g��3��a�v�����jr�t��P����,H&}I`~C�D4��'[�g.������bѤ��Z��kU5z�ۜ��t�ɐ2��d��,� _%W�8�8Գ�I�ԱI�����&+ ��&��DOzߛ|R�tt�Y��$��A������D�A[�&�zY��p���z9�1�����s<&bK!�Ҕ��3���0I�E�7��>t�؍S�������"����<|�]7���d�]g�2長�w�Vȏ�0�-��%�-��ن�� ���K�z��wQ*S���0 �iv�q�j��sf�vF�9;:�-�d��H����t�`�)c̝QN� �kv�O���N��Ʈ���h"�AT1?���^�d���C[���󟅂_a:ۙt�-F� ����h琂�x)�oB'QP'xS�3Dx1Vw���%�aP�qv���z MH��@��ތ���8	X��'��kr���A!���J,�L��8�ܼ���P,�	���F�����糖$ໍK�:\��'� �R�w��OK���8rf?�=���Hq�]?�L�u�	Ө�7��]A��\7
z�#��BǓ��{�)��=�����b)����Ȯr-��wyP��朜|3�E�J��W�����Y���_g��*�q^�D]%G4O`i��c�|����hP㈱�>a����
�`Y��l&mR�IJjv��uǭ�@��b�('ա_F�X�5�E
����NZ" �(E0K5nO�[]�7̳�8\���4�X��}�+� ɺH-��M�J�F���Zq�����Ο
�VЄ�=�V�K�Y��X�9.��;}7#�Rlr�1��Hy`	��\����,dX�t>��_���X� ���M�4�٭�|���x8Uƍ��v^���T�p���y����x﹢�y]v�*�G��Uj~l�Z\*�X�u9>m��x���Q\nse	>g�KL����	����6�7!G�t���:�T���.UA��]#�:�:�.�zF8�%��@H]����K��=�����D��, �t�=�5��B���D[���H�PF�H����j�E]/�j�Y�m`{�\��y55[����L�a�]2Z��$&�SJ��(��3L������%=
�K�$_k.�����p�e�^[���Ь1�y�ldY�\�G�20'�����2�7�p?�B�U�%F�߶���jpX��"0/O=��������8���_"�� ��B�j�GW�\w*�o�Ddߛ((KuL����-N��6�8�ۉ�<�XPgSJ�*)���JŠkq������M��8�II�(���9��#����~�^�)�6��������E*G��:"8��x�}�A�>*><�(�/!Dz��c)8��x����������C����>�)���R�rT6~?<�!d)+��1ɳI�x[��1lII��Hب\`Y��gW?~���!��ښ|f��EU��*�0~�E�����s��YmW��H�{�s�W�lˍ0׹�)Ն<�r
<��^{�SA@���CY�%��mtmrFJF5�h��S��y���HL�ˈ�1�L��qkS���ukt:#�6},}Ptޥn�,��k�-��F<�ܫ�R�^@?��E��a�7HҔ���_[���PCT#쀏�\�"��^6>�1ߊJ�@�x�h����<�s��������;%	��[�O_u�ۇC�oą�.}�G�Ր�>!�����E�U��(�pf�e��HWX=�u�}d�f� ���b����{�����Y�)!�:����1x���=�Ƣ]�^U\���G�iJ��kS��Ķ����}�Q)�^�{�(!��ĝ�/K�E�G�I�n�&��5}Q�ۭr0ʅ���-X�&�G7�~�v���ޢ,