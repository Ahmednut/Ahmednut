XlxV64EB    fa00    2b60�؞�e�v:E'�R�I�����b�S���d��8����ņ��FZ[D

���C��{T�B�+��-lI�̚ю)�IA_!՘����Ov�K���qȡ���Lkާ�̜1���g�G�I�Ğ5r7Z����DMk�,� �t�K܄У�����*��W�Q���J6q�6���?�:ÿ��cM���1�d���:�g2��/>+@)���@�ᵴ�^�V��pl���R���
^���:`E�|t@��q�~غo���\%�aǮ�6��|=/[��v��^���2�5�\x������\��p8�.ۮ���Rq�H�
���Sxх�|�b3'0���$OC���І��1<�=�/ZF��������*u��p���,�\O�x�H�PU�%��F� nz�����.5��hܻT�Ԡ�#a�%����a�AB�{X���q�9�"����ȎrJ�\��Vt�G����D;��y�)z�� W�Ը�\`@�ƌ�}��6Z�q���q��q�/ݱk%�.��
����#f�U �p9�{4��h�,3�c���]�����7����a���������8׌� !F�)��>��ڷ=D��DoM�X�_�<:%{C���yw����+��M�r���~e'L��;4�(5?+���}QPM]������zQ�@�3d�+Kl&�ȉ�P�l'���rt�,w���ym��0%V��#�L~�U�� 	3f�FO����Z�?h\ ��k%��]>=2T�b�K��٤D��m�tX�;`��oA<��T�TQ�B`��|�7���߮ )L{����J��o�R���˚�j�1Wt ������Ҟ�@�����������{�/�s�O�f�ۺXdz&�<���n���e�����.�#e�v}vܐ�܅$�G�WZ�}�b��nr����]0=+�>6h(F�Pð3;Mo�w�J��6���	��SJ%u�3�7��V�`��Pu���TL g�\�&2D!C����p�p��\c%6j�7'*M��n���CU"��K]�컣���|��N��R�Hp���5U�q\�-X��;�0����Y�eB�������Ӭܹ�)]�#|��a�Z��o�ln��er;�>�z,T()$� ��kj�W6P�]SP?meym�|-:=�	��E`���ai�.���򂖭J��C�m��ՉZKI�Ph��k�ëb����0�V~Iڭ�#䝹�-%��&�T��RvJL��:��u�j��9^���9<�:#�I���.~�_�A
[2�}�50]��s���>�t���C�Ot��ﾉ�E�p\S�>�Ĳ����\���� 1,����I��m?wM������c��x�.���=�	QG�0op\�>�wɹ�j\��z��`E�{������z�����d�)��47��?�?�R�������^��L�3�����qI��@�E�b+ ��lYJ�U��/J������l�>+k�.���N�N>;�nan��+��J'>Mc�L3�WCKLB�Bk��������^h|���W���{Z\m�Ì#L���0���)w���G���\�H^v}.nѺ��[�3�w6Q�H` ��x]�;�%0��O��u�0zY�\�^z��9��ӮLDj����W��Q�ϊ-愳���wQ,C�"�6wyK����*��L�'��ŝ<�S�U�����r�x�{R=���$b{X�3*�c�㪴ܫ����#�q�>ת���Z���V��})
꫚z��Q4Z��_���k�*�i[3���<�����c@��8?�a��)���R���cIr�-�ְG�X������׷�XXTwݥ���W� ���f � g>���]�3�[�Lƞ}���b`���m��5�ykH
	K��9b1�{�$bS�:yø*z'�^^�����ɓ](P�;D�Q��`���ݫ΢���>�^HNU����!k�X�����a��cdڪ��Lm�����O鼊��;�	��^��I�b����:�ۗ�6���Ԛ&V>�{�Y�J��K�o��Wl�w�'�r����L0�&���5�Ŗv�Z��l�X��ؤ�E��a���9�e�~���t�\�	b�G�Į<�8\��Aq��K��|w���쏥�deX94,*�k�@�8�r:�O��҄'q�q���9o��0o���?�H�1����jW%˟܂���AT`eLV���Ǆ�r��zNT�d�x7��e�*��
�.�A^�^;�&�<��0僎M#�ěj�{�X$%5��f�@��̨�1�.R������˰�Y�t�6��!���$�%��dy����<�ʻU���DF�����:��:����I~O���/�r��n�A�'P�$��A���n��A�\Q��{��W_Gۉ����&�р�B�Ls��B��4�^e�ƹ^a%o�s0�H�����d3�,>Tw7٬�ߒ��qw���#1@$���P(���~��&������I3@iĵb[,���~P�3��p*�E�W'nV��u�����󷦫�"����4�V�B��\���5-����7��Wd��o�r�S�\��BZn����PZKT�
2���p�l��T�mV���E:��A�wݮ�F{8?�҃�x�s��o�F����$�T����|f��6����=�y�E����p&jO���S�jp��1���y!�
���M��b�
+�Z��%��0͗ �CsP\�Z���t��9�DGq����,�p�p�����/C�t`�_�ז":о�lg�4dN��Y:�p��)S���8��kW��X7ڗ���T�~��kG����;-��N�G�;w���UT?���2�΂��j��D�q������rR��F*ѼD�	N��E��Y�R����q:�0_�w�qo[����К�#c��G����"�����p$b�`8��K�ս+�@<4Յ�ꈷ?!���^:?!�����gU���W@�����1���f1F�j���A@����^���N�!��TB��p�	9}�
��%+��� 9S����S �7��
���<4rC؇jQ�����?�gT�7?O�[j��#���-��=�L�Ī|H|&1BS �m=�3�i~[B�xK9���1�UZ�B�_���a�c��J]Uo{N��J�ݚ�i�Qj̏G��{��h���=�D"���=V��%���e:_c��/� ��	�ݴ���V���(�v9H4�ah'��#��b��y�b���'K	:"�ʄW
�NL�k�,��Ng �(#qH������VES��ud�ڂF�]������:�J���H�L/B��ʔ�G�gSy���`i��_��ᝄ�"��+{q�K
�V.��]�����*Ș�a6'��.$�zMD�H�C�"���ӿ��5#���[�2�ž?T)x��n_��Lt˪D�0?Ə��]!�%�/DE��if1��/���-J�.E8&��
ѵ�1��!�F��?��n� ���e��e4v_e�2�k���(fxq�ϴ��ի�P��g@-솾ߐT�̹�H��'�AL/ʒ��r?�!�!%uWˠU�i��G��/���� �r�z��Vc�Ǟ[kn���=g~��Z�
͇�{���
ZC<�����Uhօ��%c���RU�Oң��I.o�-6ߟ���	��9�:���(��2[�;�.g�FEAV
Q%�i��N#ϲ���<��,�E����bAm���t0��=�0?[fK	�3��Y`�LT4XيÚX1s0d9�RO\�{��H8%��|��I�%N���C��/K��d��#ָwz�fu$��� L9���I�p_E�Yo�X��\z�ل����{U��	��Ă�sM�o��F:��c"���[7j����d=wi��3�;7FCO�����X�PE�����Q)᭓ ����uk��d]�6��M�	���4�1W��D��B�Knn��m�P�L��c�g�t������v~TA�Y�Ewao�S�$�x�%�ek�F�|�rkRy�F��`��;b ������?�����_q}��1V�����r����6!|��b��m�).EH��L��z�,c���N{����8Q��e�M҇�5�(��ƨޅ!�a�c��x�@!����t8P�5
�cF���"�����hA�y��{��[1՗Honے�n�!{���������B�����F ���`6e~Q�*�Q�g$���M[��4����3 Z��g�=i���
��)��_fy���������#���{�m[E�A���1��<0��\I̜)D~j�CCmT�UG�����]�b�/Z�<`)��o�J?���0�_�1���t�"����[_�wvzUapKw����
�����Pvжc�!�q	�b_�&�[�N�U�4�������Pc#�,������[��+-p�����b�I?���f^�:]�_��7J��p�:�b bĝ@�W��y�k�J]��T�B��.����[q���m��^���`��	k$��m���ܟir��p��~nR��s]Bǆ�¾Ŵ�]�#7��~Șt�OȺ����'z�F�!��w����.u��wt����!AQ/�&�)_���k�k
S`#WE]x�Xv�� ���A߀6�,�s���c��[�*���� .'����iB���y�9��d1��#�ٳc�t�&�*R�"?����Ũ���= }��'��$�����f#��x�r��[?s��>���Qi�%z�c&���b4��Z�S6A
.��Lfb{��YW$a�ZpԖ��l�j<���Q����K|n�=�	)�5��\�+V�-��
=������1���@�Ih~�U�s�˗�����|t��V��4.�p<(vA2���8<�y[d��?���.ލk�����	��H���R�8��ma���l?���3;}�	_�U�kS=�b�c^ɬp����t$ F�����_Ρ��w563t�CGG�$���G,\*���6D��m	�Q���}>j�ֶܻ����/o���I�5�V�|���u����Z��|��*N�yڐ
��.�5�γ�&;sf���b8۱*$�>>^���x�6F�x��FP�Ќ�Y��p�۴$�e�˒�6���?D�H&�e�>8����C� ��R��5��<3�c�����G�`"�~Ehm�y�8l�����g�D�7	_-ڊ`;툛s�!K�uC7���0 �Ԩ���&+{�3w����?(+�Ne����N~j9��a�-��:@i+�������H�E�5E���|����! D���C�R�}���+�AH��O	pl�"��V��`o���՛.�*�Q��4ka�#$��P��H"`�#��s�=B^�)~�bN�QBJ��;��뇇]I=�͎Y��&�viK�t4,斧b��_+�䃘��Q�yб�X�if�}Ї(�����y��Ή�����4��3m>�&8{� �2�V:. ߽�g�Z�_ZPWN� ���v8����P����E��3�mTJ��%]sv]
��;w�m�<N5Ɵ�R6R�������7Xs��ZR:o���Q�kT��%6�/hS�vj+a��y�F�Y�h��(�xB��a;N�<*�Qn�h5$��"Z�n6
��m���1�SN(׉s�P�\���;6tqEl�i��:�j����w��Q��g�/��g��U��ɷ�ʞ��R�]�q��,�iɎ�>���g��S��9(�@�%m������2o��[��7vo`��:VZu��2˘�&���>�xL��� 2R_8P��7�V�+�W#l����/H-�}-k՗A���W���Q�5F� ōM[a|��!��mè���o�ܿ9�'4��y���C&�iV~ѯ>!N��6�0�׉����2n���kU�h;��r'߷�ٛP���xuw�* �&�>2�7`�ҽ��Z���Fc����>�K����sqP1�5#�k�<�ۮ��^j�
��Zӿ�3U8mv�W"MމIը^w�0c�^�	0�s���쨯�y�#W��ħ��H�]E+F�f������G�B�wh���R�o���Rq��:�	����`���ВՀ%��O�9��S�;����0���X���Գ�c�9J/��a�L�C 8�W4�,/%�Zy��f�W�F�1��h>�lE�����\P;�Ѧ� W���D+-l�2?˷u�*�*�>�ŧ�ٿIL�PC���"����q�bF�𧑏YmI)t� b��G�;����ȰB����|Գ�1�gwA;c3N��m`M�s���Ԇ����M	\�����m�	��aA@�![&
��Q��^�G ��7)Q�ؑ0��5��]3�P}��؎���5a.^�Ҹ���b�e�m��f�PeX�
�o��,��:b��2����JH�o_$�WX.�!+o{�eo�89obF�^��+ �G��s����p� o����$�~�Dg@ĩM�ٻ�;l��~���N@��t�τ��u�gypb�(*{�!4=�5�;];�#�ۋ�B����H����"�F�ߩ*(n�ZfwMSB�R�X֏!���d2|t�v�%0ݻV"]���_q�+^B��p��8t���;q����/��A�i�ޚ{�w�yY�n�	������o~L��%;�KZԨ�ڤX0�AV�(E.J.��h�e�\�M"�xR��3�Y�c��KL��2ʸ��	��z%���^6BAw�Ofwnp?no������s�u�
�R�->^/rT�	�F�2n�&��m~��� xs�v�mh"���u�����h
\�*k��a�3�d6	Z�Z���k�m����*r�������Hٙxs�
˦�#=��Si��M-��u�}��>��}��i����� E��AZ'�}��ʱ<�nEc���y�;���̻���TP��L+gD�	R{�]}
�Z`~�}y��mɏ[�(�.�*Mq޵shbE�j}b�t��$����2��s�Z,����r��!��A`=
۟�W�e�%�}�ɸ{`RqO�����b��F�r��+",m%ײ؜��Au�:d���I�L��h��w��Y";���
�
����|W�7�/�T|��b��v�����\���c o��-gaP㌩YW��d�=y������x�*d ]��=FɽZު�

�Q�m�P@H7���C�����
]�"N��0��y-��:hH���u!1[�EC�~Jr�G{�'�jK�z�e�֊0� 6��}1�E�_pJ��O�`��0�ߘ�e�l����{_�٦0JF\]�
 ���x\_����Qj˵������L+Y��:x�k�@S�����xm��t�#VU���d��1X���#�zڂk�~?kYH���`�3޽~�1׈V�|�Dv��=���eȺ����}'-7�+0��Ţ�|��:�t�!�(Za�Y(L�rӶ��Ѱ�@}/�#j�}y��-u{,Ϳ�S�]zUΈB�O܏�����#���g"���b����2,泘	�4�����G�:c�;��d���tԃ�L%��-ӿ����鄯���8C���h�Х ���Js��弟<��j�����"�M<h�RW�S�g�7�����E�����B�Y8�IzsI�:�A����z����9�`��Gg��C>�JڎЛ7&���%�:M����ֿ�3h�H�*]���ܶ�^�Ґ�`/x��*��vJj�����7�\�Ւ�1N�������Fk�J�����d�r���N<���z�M��Sc�I|�<����>۞��^���}mP��B��s��t�L��Cѕx�ܡ��<$*�h�l�/�?<�Ʌ�Yk�
���w�<>6��y��m-���\�����U$����E�n$:8� ��4�A�$�-D��G*��x9w�.\EբE�5΀�5�o=(���{�GE�p��[Yc޻�vO�Pm���*i�ρJ�~12ʮ�ɜ�v�힟є��5K��!u�3͙%�d���OM����#-��<�O��m
���&�O�T���K�y�-kh��P��}�C��$�P��33��mF��*y,smq�*�%�[�O��V�y� �8�ᑘjX��r6��U6.�%&0�Gx˙'nN�M/��5������]��gݏ�@��"�w�"���ƍ���V[�c5�B�,o�P�#DEwx�kYBPW�����(	h˦7L�ӓ��w���Y?)�x�ea#�ή��f�B\$�E�����i
�g�)�#�f����G������j\���}�*�o��(},q�<}A}v��ݱ�����A�9��_�4�Bv٢j�����CzX��0h�E�����cv	@$�t���:�\�����TT)���R&��!�����xb�	-t�o�gO���h2	�;W3��C�qb����*���9.�bl��@>��k쵠0�3�;��O�h�2��b��	r�N�-�9����8�t`lͼ��q��Y!=6]˩��'�I0P�7 ��<LPu�/⣠)��\W8t�CO���u(��4z4O,�^R'�Ғd���%�W��@#���Ԍ�x�����e�R���FV�y6!��B���@�F;�%(E2<�+6�I���3�r�u۞��t�ГY�dS����'J,u���5�Xt(�F��=��?,�N���P��s�oa
���e�H��(�����u5�^h����TMyY�o���T�WI���nǞ��S�<����h-��8����;����9��5<%l�>��Jۼ�0����1�J�p@�!\��B���	��uc�2F�t������FR��V���!�yǴ5��n�ݘ3<D��+�t�(��I���W&��s⸂ȡ+��T[�p�.#oM�J{iÉ8f��@�2��>cj؍K/�6�8.1�53����?�˓�^Ya�Q�Ϯ�y��K���e��&^_��ݾ��x���O�b�T3�5�O?�ʋ[�H$�I�Z����ǣ��d+�`�\}x;���r�.v"�Ҭ��W�&y�n�*��U��c�n� ����3����ո���r���n���Q�xX'����w�9֐ĥ^�&��" ��������d�1;�{���,M�v�y�?�GfMG��4���,�U>��ȱ��#H��L1-~�OKނ>[UQ��25*�yι�9�H'��4��_�˱�mq/�Q��!	iZiޯ����S8� ��!7��m���p�U��(���:������8���y��~C%q	z�+j*|e����Zǰ��刕Jt`L�}>��L�һ��EŔ������]⏷B�%MX,lF��Oo��<m�vFڠuU��\E�hR�(F셂�:�ՔTF�M�=n�`8�0J��0H��UwaA
���^~�6����R�!���Ԍ{`����]9T<a�h�R\*VP���
��20!�I���5)�P�͏��^6���ܿ=��twm|��?Y�y�'���9�O��3D��Nd���6C�̏u�B�o�@��,�Œ�6wջsPR)�In�X�Ah� Z���-�.hv���l��B���唘I�aG a+Yu
^�3�Ɇ�a�I��ჳzȤA,��
d�*2�Zi�D��vh�$��W����նsZ�� ��%a�u�}Rx�*>���#g[7ZBF�O���B���y0�$�m����	�g3����T�9��.�/o�P�u�6���֔	[ƃa��b v��r�ӄ3'Ɣ�l��%|�8N{P��H}!�Dp��cwsX4S4n��b����&!�������v�uU,)ZVn�͍X����R��u�-��]�

Qf��%"�aE����+����4$%&�e,���ik�խ��w�r�s1PL�S��Ǳ��D��}�Pyz�s�^1)/D��#�86�����������Q�&��Ē|M�:+�6=��ME��mqO�z���ܢ�7��7���xn����4d�}��2����J7ck�Ǜ�,^������~��"�T���4�Dh"h���y?6!��62ףf���$�@w9��h�5~o��է����<�q1���*�}p|k�O{||�Eڔ�%��p�4�&&��	ser�5_\�D�J)��~|Č^�=�0ô��A^S�j�6����H��T9�N���w�]�-�2��0v+"w[�E���\�n�k�Gl��aD(�5�0����Ik����u�z�zĭU�� �P�"�=BFlc�냹p�9N�(��A@�{�!cf �*�#)ڣ8^U��ce�ٵ�7������rK�v�0��俔��@�5��CI�P�HF���~uٙi��G��{��D����_-|î��[LMko���xl�LXȔ{�|���Axĺɲ@�fi3��w�@Y~��ϣ"�rP*d�0`m�m�@�7�<�c:�����h�C�R��J�q���/�d�]G�>6p���B6̅���8"#'~�V⻋:�����3s�������$�c��Că�=��SM�>Br	І�BLz)�xSn��$��Q{�E�.�>nYy̂�C��Z�Sc�ʎ��x��|��"��w���'9V9~�ag�6O�}_�*�A��oc��m����K�� u�d����t�<��W`�4<���3��5�a�y�t�=�r��4j���h��B���V�h�0�� w�ȗ���wh6�%�Ů�*%�>²ƁS ږt\�H˔����#@�����Z�BK��������7sN	�ôj���
�:k���ur��TO������
,�C/a�g�Ύ �����A֦F����������J u���^������Τ�"�NhU4�ڲOQX�-�z�r���$�!����ʭ&�^�cT���8��V�V�ӱr�X	;{����������. _::��1n�W�T�����s��'��~Ѱ��^{E�Jw�Bz.XlxV64EB    fa00    2810�L!�pÓ3����O���꓂���tjҌ0Yvۄ�pfH̹�c���+���w�H�}4w��o��/j0~����ӕ�T�>pN�cq �
HgH~�6M�C�P	�`�)'���,��HҜ�	0��j�C|�{ %��@#��0�jv �`3����8X;���H8��81��2�� ��",]��Pd,�F(��$�8�j��-�ݣ�]1��$Ym�Π삆�X- 0M@�ꀃ;sw��z�JzCh�&;��	郁d�C�z@����qG�y�2�2m��]�����n�r�ݓ�3m4:�|nX�gq��Ř�w�� ���8�<X�z-:���Vt�x&�[�����K�<�����V��$��vE���G�I��c\at����A�޺x&��o)o��\���d�$p�����%ޡ��i=��#Z6)ƙ�v<7w[)��e��*/�ʠmO%�_�ʪz��s��%DU�C�Tv���^��I��#,?!=N�]�Y��d���cDB|�Xz�S`�Ŭmr987cF���y<A@Fv�|0��/��k�22R�%u-l�e�Y�z޺q�b0B�JkQw�ؗ m�C���L��v9�n"��-"ܱ\[�@���s8������`I%^!J��b Wх�30��!%e�[#/
��R&��J�0��T6� 0�&`��r�[���s/G�T*�*5z��n�խkwx�o�|��k�UϯG��DIj. ���3Ғw����!]=�0rg�[RǺ�؂��ӑfJ�r��r)�@?���2|s(h:ip�G���.� j�RW����	�����:0�=�12���4��Y"�e"5���5��x
�C����A�a=`������'9:�m�|T�XM]��B!|�����t:>:5#>��3Ԋ�9���D$y��3�a�|_�V������5U?G8�{��� x�K4�r>�)����0���J��k6y�ǃ�̂�A�-�3�s7�=��q[�� 3��/��Pi�� l��o������+��2�$O�A0��F�b�f;3/	�{;�#��R��P���#���0�v��I�|�VR�@	���x��d7{y����GZ�^�#��gVBlO/�v�`2���-���R�RE�16&���r����҂l��[+��������K�$1�0U�3aQݙ���\4����π X-�B*?&Lcӆ,[�������&hЩHچ�%?&�14u���9�zTj]�R?��[�%D>�S �G�G�I�PkyUCBe�Ce�&̋]��g��p��T����T(�� ]f�04�?C5I�J͡��V��G���v�"��
�^�����	�0�F^�q�k�J���x���B9Uy�l��֠y�ٴ"����̈́�^|*��;��]0B�\���a��P~��i��8�F�tlS��*a���|�Ұ��3���h���Pz�Y���d��+&��$���d]�Iy��f��oC���`V��pI{�nU
z��Y�c8�`Fd9	[3�Ka�Zy h��QP3��l�'�U�y�#`^��1'zr�|w.��ߌ�n�Tt��gS��ّ�;���sX`�͇��G�t�Jʕ�x�N�"��[���ٲ��Cƌ3>^��Yr��s�ӈ��~,1��o�Lߣa�~6E@ϕ�ꢂ�����L�(Gv#���ڡ�	�ڱxv���C=�� ���ū��x�Av8���T<�ֻ��l�S�Y71[�@!���C~-��Á�\J�ٌb��S�x���X){*D���/�â������!�М`4�U�����E�fHkQx����ym�	�ީ�<l;LE_Id�_q-� Bda�9�Q���G�x��C�V^�:B�:r ����H�і�`Eb�aZ��̎A�p�xZ Nq�d߻�\�l�gޞ=u}�qmՕd����������G��g�t�5��"	��wV��Y�M�LVf2��0?�Ep_)�v&}^�6�۱ �+;F�&L85K��w>R���U
�Jh�����5;7���4ϼ^Z�R?4�a~��`��n�?Z�Q8j�SJǛ�������C��MG�`�U�@���н�,���+X�i�+t?����,a��nԎ��qfs� ú�q�>Mz���*m>�|d�+װ* �yNzd�p8��nb3�
�:qb�{�IO��h���a��nI�~�r��m�5�`�[ڀn���?�Ich}Uu(���N��Ew�	�<�G��xJ�( �R->��_��9���Ώ͑5%|�G�_�(gf��7�2d�N?,`ȧRd�����z�DE��%�EZUE"���Y�n�UEJ�6��cF����ļQ��sa�8���V�UJ���*�.3�h�M�eu�[(�ަ�*���G�D�3s#��"yF|��G�Z�t����1�A@C���%��]=��1%$[di{,�ԙ�T'����r��C����Pz�۫��;�)Wo��*��.�/�ų�V�l�_?@0b^�0��׻Z�~������E�Ɇ���0�O��t��ϐ!�j�#�%2W�����.J;g�>��QZC�ڮ�����6kZ�`�ZwŹ�,�lE�)��#3��(ư�D�j���� �������sm(S�[1�ڨωģv�G���J�v�
�ȫ=\[��_N�G�S��yV.��bc,�3�h�,_�D�1�9����϶8vfZ�JT+ID��r��d|��ULN� Uu�_��o��8W�2z�ɫ�t���{]s��g��:Z�00>j < �c�	4h�����A���@$H8����}���ģR\�5��$�E~a���~��q�s��ݢ�W5��4���X���6P-��������L�Q�7ޛ��ywv�-@�Xk�{8����!�u��a"�?h��j^~$�Y�<OmLN���+[_��j9нhS ���y�,�D��VX2�^��.g���(*;Л�*��i�i;��ݚ{�G5���DV� ���y>tM��h��S��U���~ld���R�-.݄�7�]xj?V��=� ~�ے���[�����M-�a� �7=RG�<�$�֘:�h�Z*0�z�!T�ϓެ-:nCG���[/�����״�{�-��gN�����u��n���F��0!4ʝ�f��jav���M���k������� z�M#���O#�.Ȑ�=����1��� �iWӅ�������F� �i4�l4�WC�≳l�ZxD�^\�� _���g�ZŘ
�τ+U�f����BK�q�[��j���t:&�J��[ȍM����;�f"����{Cj-aA�P2�>�=۲wIѨ�Hpy��8g�1�2Ok�{��*�F�'/�����?dw�*�(�-�p�'H��穹��45��8.i��]�O����A��_;.g(�R���)57j���L���XŻ{1���c�zhM`�Q2�λ-rb�k"u[+��wޗ���@[<�C�&��6�=����������r� p�Wx֬Rge�_�-5=c���\	�e�y���3��FK�k�xW�S��B��&�� HS�rO�A�="qK<���Қ\��ܣZqm���ݒ@��[X��S��[m�j2��O3\������p��[�٤�m~ ��yq겂s:�#[�%���xgF��N�e�Z�*�9���9���&F�(r5vlP
~�� �uj��a��M�f��F��]� Rր��.���ϼъ� �/dH`��C6l/�ug�bWok����H1Wm'��<�f$a�x=,;���C���#���Mb�:/��v�jvV�bP=?�r�Y�1���u�dK�T7p��	�k3&Vڮ4�!���8���K4��|6�F���t}O,�U��۫Q���.��ڠ���׼qm<�|lv[�Rh&��
��#HN/ĺٔ⻰���*%�U.Kh�@XO����{B�f�I�~����C�#D'��0���G꾤�הJt���B����"0tP;AF�z�c�a�oI��O��i��=�ϫ��`����p]o_c��{V����L�k�b�R�q��$fʹwʥ��)�_򱬽񴌢ŝ^2&`Z�a4����)_3��qEG)"nd���I��s��}��qC��L�;ܞjZ���o�~�T:�q��S����$<�?W��	���e6�_W%���6g�3&ɣ$X�2
����I�a����qy�F>�-4[��6��obc�6�z�ߘN�d�����wg�
�Q0O%%�wz{�1\~�Ě�J?I\�k(gӋ�e��!`��
'ã�����?���6�sZ[�Z=�BC� Y弡��a@nˉ�ۚV'�@8���։pL���X�8�)|���b�-\]O�s��.� �=�����1T�>�f��F�ITs�GQ�/��E�+$K��tR+f
�E65E�Tk�]���G��@ܬ�y�pi�37�Շb����VD����8�x�Z���2jx�%���o�l��rY� �rwϭs�z�ܪ�j1��w�
�'E�_�N2â(üS2���r:e���Чƶ���<��G�|�H<k�ўD��J*8��1v�.ڰa�W���$
g����|\�/�h�z��èEx��֍!h�����e��4r���j[js���&�D��������t?�x��PD�p&j�wN!nTV(���vx0ipӶV>��d���Ն����)1�_�w��زT	 �z�h�*��<fZKFg�h��ѻ)��1p�4�i�Ħ6L�:�OWY�,|kJ�o}���l���@�&P쒼��@�,������&�M�"Q$a��~��1I�h����Q��]-?�1�af��-�;5)�i�����Y��~��>u��j�)v!�:�o����Ou���;{~�!���4#y�D?�뚚�%�х�����MoJ�6#|���.�r��p������h₴s�,��l[���^2�O�,��+����{%\5Ó��o�"A*#o��z]�j��F(6����d��ct,���e�;�jV#aᬉ������a��w�X�NXY���mh��V/�ĵn�x�]�}�yb�Ph@��3\�8��m(�\jW���f�[�{��9T�+.�4]h*�am~v?r���6\RBi���[��e�H��.����\U�Z��]�߂��.5�l�=�%zz��	pG�KkD�6��V�����C�04���Tq��C�t2��{�%�
�����/7���@���3����>�o3c��f�Zc�B��>i�o��v�VtmF3�oL�3���T��u�C��x@��6��%�|��-`�씨_�{9#5O l�aU	;g����s�S������	=�<aae|�����5�f]4"�@¨����UDj�DN�F����C9���>h"x|G����r��:��?�rv͍�ܻ˟;�f��Gcu����1g	���t���:�ҒIwO��ync�9Ek0P�it}�,U�R��2(D܏������\�݅�5�7�q5�s�2Z	��|��R�o-#��mB�^3z�&��[��vX��Ę������&֛V�tj6�8����e`ԁ�+�g�ސ���*{'�(��Js]�}zh ����#l2��>g�rv����U#R�pU�*YG�aSJ�]QJ���"0�p�&���S"��<�T���@��"�`V�W�c@ͮ0���kJmA�XK�d˃�� ��I�d�my�hj@������2�h����G�+/��5D�b�3O�����VME5�~)
�*nUt�����-�ڋ5� �{ªc��*��r�7����V%S���$��w��
L������0�+/��J�ۭ�)r`^E��Qݰ�����C	E���Z����7���� ]BVQ�j? \�f]?��_]0� ��.E��ȭ~�F�<nL�?v ����=�~�{��Ub��v2३�[)P||Y�6oK��7�n~QS�yH[�ݐs	YID��b0�C�C$��f�j��#Y�;f�D�ӗ-�LC��<� r7�������g�)���y�[dZdk��%�Q�6ܜ|O��_8��k<�����)�b�G�3��'�]hq�&ss�-9�-vi�X��o+\U�F�)*�'d�+���kݮ��s�F�s{"D��V��&+_�e�9�C���Xaa<���3�_1�vEK,�	�)�������Ri����Q����X4Օ�Jf?^�֬�ʂ�<�6�d՜}'�XMe�$@�r�3B��V>*���Պ��:���]$3�Ժ��jzq�eʧ�D����ۯ&l@�C8([p{��~U���c�+�`ܫ�C��$n���彚IO���TIom7o>��;�&�� `���5�	1��5`�p�d�e���W�I Ek �5��N�����+O@�0�H.���O� ��P�.rk4`i��t���o��[�J)%��R�KxF�š$G�+�i�����.1��?:d'���t{5��&�c3�g��ߤvj�(�Jѵķ���
N'�"��p��ID��R�(-��P*T����]ϋ�Q0���{�5�/�uW|͟N|���3��*�sx���p_���a9���VEE�C�k�3i�����8��e��V�"&����S��t�H�R��R� �N��-a�!x����`�d6���b�;1��l����op~�¢1L��bcӖɕa�M�S@��`<�6u�LҺ��1���O��#��N؞��w�s���#�Г::Ę���]���D+n憭@��־X<qe9i����D�߯4���V�58D�������b$;B����������k�-�T �fg���J����I�XX��_٥LH�A���dD��L�;`���+��`�%�ZJnb��;�T��Y���&���nw�<����lT�a@OmdsY`�2�N�޸B��^�gu���|˗gj���r_z�у7yц_,ڕ�Qh�Gf��ٌN/�q��_�nC��^}��R�d���|�m'J��T�t@U��LC�´1!d���2f���Jg3�s4����h �gh��g�X0ύ�s�2�f^n�
��������"�w����fբ���"]t��o�;Z���0�!���sΗ��%�qѻE�劥���S[�4B0����)yQ�È��I1zD�ͅ��?'� ��Plp��)u���v��#�X�du��DC�Z�D�l���՞�\o�֤��8�-<в����L5���{s�Āݣ&�"�M�h= -���9�Ę�o'�w�	!���v�����dl����_�=
W\��g�a��mE;e��JjIV�k�Q�>�76��0O;&b𹧘b�10(�(3J�u�d�~_ɐ? ���m���j�F����%���~6��q�a`������/ �Q.�)늓{ߩ'��}�J�ya~z���c��w�|au;���J���Ls�ca|�[�1=.�rn�����&ro�Ń�I��mX˓�'�`$�L�I����H�J��*���pb27)E��g��u���d�خ�LqB�P�	Ɂ=0���Y��c�Z�4�Ѣ�
8<+�M��j��b$�e���hT �aoX8NVZCZ\ �����B	��:��3.�n���"�+�~�R�
��^�H�\��~�F���5d��ߎ���ҙ�M�r��Q$���� ��(����s��p����s}#ŷ��r�sg �!47x��@�a��8S!K��<�/��m�s_�5*�(I�2I!/�U�,~^�ȯ`.X��*52wy��.�m�nŕ�G*���jm�g/p�5?o5|�}c�l�]�vzV�p��Xw�i6�Ԇ�+�9�V�p�F���e�g!M�N- ��6����B�ɍԅ_^B�2��n#[b�������t�]TY��h����꣢_��������uc�okNP�a��h�s}�<n�(�I�J+��}7jg�b�)����mk7�|5����Rc��O�t���$T��25����$ɡ4B]�GwU�������'���R���E|�g�vI�Q���Y]� ��@yRv$�h����o0����a��ƜWN:|�<����1?�y4.����t�0ły����tu;��}m99N2����h��B�s��{�u���I[l7�t�ȥ:�V����O,·}��\�Ը�G-����k�O�-��m��ӄڧ���M��m	��^=q�)�Y�ӉTO�7C3pk��U�NR���"���2��ߝ[ˌ6;�I�1#��b�ґ�^ok��A6��n��w�����m?eՉ}1��e�s�nΪ�,���+����-O��58Z�v���[I�e�?7g��٥^��1��*���&��m��J�ǎ�ɟ��e6V��+��q�!��wvYk�@�v��WKJ�Ŵ݁�*z�Cdǂ��8�SOb�{<I�>jԾw����-��;0�+��n�Z����P�|�t�VW���ߢ�n$��M[D��ă%7�_Ю	���c?]�xJ�SJ_f�w�M7���vY���et�Z�d``8�h'��u��&�Q�+J��2s��0�^k!Ai��Q� �@��8�������!?��Iޚ���uYZ���#��2;� ���+Wz����Hc�R���j[�oS�t���k�v��~�
�K����M7cĊ\�89��)��Ex�"nD����q���P�tǔׄ7��5r���$�*��}�/['VĽ倣Z�>�#�H��hj2��ˠ���G7�{Hg�*���d���+�<���@N�/po��0��H�-���)ȍ"��]?�S`��.H�j��v���r���w�B?�U�l��!Ɂ��Ea�:a𙸂<�Y���y�ӹ��.Ԥ��n������d~u[�M��rj�č1�����\��$�|����uƈ	����q�+��I�B�lG3��2��os�b���pq�uN�ئ�4?C���*ƙ�~��G�D�nt˼��1U����z����X�-���X��%��9���٭�sg�X�8�fk�9�/7�؀���.0z�0bN㋞�F�%K(1���'R��R%�Yf�Eb�{#r��'o�qQ�l.�}�#�W�yε �rU�9V��w��n�������zv�����t��oǈR`�%�Ɋ�0��e9r�{�4||Xܦ�����޻�8�D^_�b��3��jI�!���O�d�w#��%B�cE����0�7x�	���_�S����-�ov��\�UM�F��v���WE��Y`R%�Q_,;�5  7�S�H�}��8%��\��h��%�U�FdNt/��N�'�����wxűI��^o2=O��T��M��*����0�[� X�q�Z0�_���n�&�ܖ��s>-'��	�K;�f&�H����Z�s%�`�r����a�)��y�tHU0�-$/?LևY�KK�i����b��v<�$�-��	�
�t��`}a�<�M�l���!Wb����H�e�w�Q��C	��1�(h��mc��sgI>f� �+)nW��G@��F��X>F��Q��%����A��BWi�5m�BVa�`IНL*N��I�U�x��R�v �Qc9��)ڱ��07�(��o,��j}��H`eP�O1e��T�5��+��`i���z�+yOR�z!��ux��e�R0FS#JףakK��cfG��*��Ϋt�gV���f�I��h�[��7��I��	��d�KnR-5��ilK�%��U4oM'��/˅�)PE�O��6������g��6��r��M�9V=����2�n"��ukE7!�ck|��ǵf|c#�̜�Q�/�: .�|�>�J	�bC�˽���,_��؛'bO�w�S����l�#����/o_� ="bSQ�[�t�iDe�qZ��A�d�2q~�C�m=��#����Eކ���Y���w%�ÅM^�t��W����n]@��0
��Ȭ=h���@��U��N���i--�6@*��_�'����fWO�oY���64��$��=�y^Lb#R��j;[wܢ�?��%��K�WXlxV64EB    3639     8d0=~ج�4���� ��}h(���2�ȿ&��+�R�_̛g�Q��cQM]`�x�����>�An7�{}`~&,��j+Ŵ[��Qj�$��p\)�u��}=��̵G2 hս��e��u�M%�y���t�+�O&���C�}��㝎�4����L��b_ckԍ����08x��Z��kc�I�������N�|����TV0���$�9Lv,Y���˴��+��7�ЙT��ip6��%A�:wi�FC�F҃�v�y�&��ɶo�s���5y�,�e�p ��΅���@� ���zg y�����?h��J��=�-����������8t十b#ɗ-t���+��+1�0�֛R�����
�'��Dic'��>�L^nG{�l����>�6�9�Y0W�9/�X܂��5�a6F�K]�)|R�݇S�Z7Oh@Q��� ��Y~S/�2M�{����L�th����`a�v�hZ �G�;���C��o����-]@�y��|m����)<�c��^�9�ͤhj�k@����wW�Ss"���JL/F��43�1���͇n�UV^���+s�)Y2���}ɩ}�N�g��3˕a��;}����+�>_d�#]��w�1ꎺb塵=�<�\g�3@��O偅Wr굛k��\(���؞����UA&��5�M��v�Ұ���D;w@BlB}�P.� ��ܙM<�4�f{�� �l3���	�K��/��5��]�Hrڼ��@{L��+�3��b]R�f���ס8�,*ǖ��orR�kv��Upn�@�zi�Kt�4�3���Y.�3�n	�����u�ɇ��P��{���Ȃ�C��B���J��t�`S͓���'1%��R�S�C���tn,Z�1��B����8��X���c����eN��?8�oG}� �5ׇ̗Q������-��2;Rޤ����Ӥ���vK�.d�*ǜ7���VH@�.�O�6ξ$SA�a�Rk������_��q��S��ة�fVQPQm��*=ʃ��+o�f~�.�����xF� Ж�}�}IX1x9AD>lB:�K��oՀ��5[
|�
�fCy'q�o?E�)���^Z��X��V���c>�u�0"L>��K�2(�!yk�@�ug��G���o@��~����u�+��ΛѦ�^��h�`�d��	�@�t]+��ĕ�c^�3箱������&Gjs;��/s�F���g��M�U�[>��X�*I�F�ޔ�%Sx�
�pj�̱�s��4����Q[d1�}�0��}^]��ۋ�o��qCв�/���5@�i ɠ�4��v&��h�Q�8� K���yS��7�GXzD������)�M� 
�Oȳ��'ih���%o�rְ��9�T�ep�{]Hn&�0q <��hU��Q"�R�3־�mk�����	g'�ر�Ќ֠_�*y����ͦ��h_ӊ�\��>��Q0��Q�I%D9�i{�e���
��۲q��z�K���c�.!?�5����T.��v�KX"�g�o�B;�]��{�h���TÐ�2{,!�lE��QP�%�J�tʀ��x����U0��P�B7ty��L��!�(� כ1�2x��P�^�@xS�o�������z�E10�ӐZU�Ԛ�%�G��w��(G�e��X��kmL�>N>>��؉�a�$2����m3���V/��W�O���^�V+S�_܄m+��K�sE��Z!�6���U:\���Q�Z�r�=\mA�)��Y��l��Pk �> ��:��b~�Y�VrZ��y?�U1�'-�R:��<�߭����\u�����)tXR�A�bx4Oc�9�y;���n2��&_H�)�.�[�&U�kiN������|B"u��H=��S�M9l�� ���r�#�D�6�D�N`��L[���GQ�A��ˣ��F����I��-+���3ut�V7~��oN�) ��(�4���J��BY�G95TW"�!ߵ�?���
�^��t�R�}1�1
7�_��������y����Ca���	8�.���^�c���谅?�$�vkp�;Ͱ��4R�����N�"�me���..g��/��|�_)�DrSw���j|7Z�`�;�j�g:�\ڐn!a��S�d�U��[��V���4�I�E'=�7��b��̇�;Ph�N�	�X�'B�R4����Hb���sV��~�]�o��!
�oYuM�E@���f�����!R7j�hR�*F&P�(�q