XlxV64EB    fa00    2dd0@RC �?d5ކW�j�x�ZF9�z��(/�i܂5H�&[�jm��5�K�L��͟��F�7,��G�F�}�H�bB;�}_}x�i������.ţڈ���%�ۂ[����X����j0�2[�3)z�,��e���IgJ��L����޷���x5��H������ׁ��%�HP�s����m@/'Q��\��(��X�+2��^��@wc�2l��Ŭ�ۍ`��6�R�mZ���j�y��D45�����J�z~¹��� ޓ|�n	)���M��J�<����(���S��#yOƴ^)��|���կ�
�T;S1��R�g�1�����\�$�#c!H���<��V� a��p=9c�	�#��h�^ݞC�O��h3AѫLE��|�K��?�O)^���I�\�-4.�&��~{�\?�:B�'c��H��,�?&�-���z,�x�
�l�qϣw�n%Ic3�Yǧ1�3c�sN>�j�d�~ƨ������+�vAm.�H�n3�ھ�LV�n1�ݽ����OH�G�i�\�7�0Ff g�������S�=s�mkJK�g����&�&
W�pB4zG�o�H�2��f#�SAZx(,�+X0�l �/H�iW4[��MZ=@����|����v'�6s;�_Qm���n/C�9��1Ǧ<��y�����`>0���7����,TfGۼ0$���T񖼿�/��3�����jg�����/�)51���b�p��-픋H�����S,�� Ic��O��E����Z 0��:6yd�/^%P�E�w�X��h{x���G���z�:�P[|�?�bbYI���"�#a�f�IS�[�3$�_�d�B)��hߧQ`��5ՅH�kYg\(��t�pևM9Mg���.߀(�0�qϢ�z���`�#��(?)h>��.��i��ipҺ
YI�Aj2/]�*�q?楧r ����y�嶺[ŕN����N��'?`�|}��6����6<�&F ��#�|�y�H0f䓴�M��N�� [�0u�G	�ꝓhC��U�ᛎ�jS�Q~M�mYӠH�Z��Z�� )��_�Ҵ��*ԿK~3c�=����<����~<p��±$c���!��ͽB�{?�~ս]��H}6{餪>$��L����Ա�0 [����0>�!4p%�N���aT8j�/�to�f:��J�r@�3�T!�RΥ4ʁ>����!��'�p������y��D��J������1�O���Uz�y�9�C�y�.Z?���U�K<=$�����ʝb?ڇ;N�SqV_��4땽���v�,�|���0�N�OEmA�� �A��+����ַ��Hd�"�Aꭍ�gt�96�%D�P组e�h�e����q��)�\V{�*�� /��������' )d�{+� �X�-N��u@�e#�|��6m /w�w*E�t�
:���xr�^P	Z�f~{�aSZ7�umzo���l���7�������8]RQ��%k�ڪ�慿~�'��-��3n�Ri�ds�b���h�n N�,O����I�O�H���"�-����]��v�p�א ����u�G��}X�@����4K1w�^����:��3�H��?p�~�#�H%��3<���ݖ�3<�~Byj:���[z�Od�����ԇ�A:�K/�lI=3f�0T��6z��2I��pP��6JN�D���CaY
5�a����_���$�mW T^�%�pK����T��__yX�:,�*WWf:�J21��-�j!Z�*������Re��$@(et�Ц��M��-��ᇾ���+2�uFy}��?z�8�!q\7�J�T|\���u#8u8N���7�i+����W��y�?���@k��C������p�s��3����E Mx�Hw�	E����	�*��.zx�������|�*#�if�s�da&2�5}��'�]��͛�G2�E ����鳞�9.��3��&vn)� �3
�h0m�s�r��5�\�?�,u��d��Qh}��ҿ�#~�E%��O��|�̼�>ru��W8�G�H��C����s�ړ���.�n"@0�g�C;E��-�L���5	��h�yC��$e���4E���X��-Kȥ�D�Rt�1B_~�z}���4@�p�����DF��E���~|,��Qf"�?/0�ji���a�~�p�q=�8D|�E���w|�	e=K��#rv��^m9὿����m�\�nb��|<�d�1�7��Iڏ�Yfiֺ:�RC�8��x|�OW����L5�N&٢Kt r&Mp)tI��ڳ[�zX�< �<�#CI�oP��&�LR�O�;5�jݟq*P�������k�ɨ#g��UNBt�6C_����I~��D��#rZQ8��yM�_��)`��Ѣm������CNn ��/��+�3~���u@!C5���	ٓW�4���M������0�6 �Yv�f�$L�?�s+��T\lY������a,�>�gZ< Y��`�p�H!��hM���%z�XčҬFo_]|@C�f����G�~�tC��M�YXU62�2�{a|����Qa't�O-z��\���L+��_�{��)�DNAoh�^-�z����vb�CT���BS-�Ss_RkBn���%(%�L��8o��hr��4��d�\6���(RO!P��[�rߑ�A�Z&��n��?�*� .��!�Ӽ+�D�g� ��w�i�;u�l � AP����8K�����ou��T���u�0� yRٓ���a\�����u�h�l�e�үQ���zӗ2�#�*�l���7Hcٮ݋rn��֣�c�~ٷ�L�[��@IHY$Co�	B��U��������k�#V'O%S���%�f=��zn*CoHG�B"���`�n�xCrND�c��������F��J�	H�O�>Pe�y9O����6[����{�cyO����`v�3�nڌ]�G�B�N:N߀R��š�X�!@���$��NE$�O# 5eO;�_F��4� �9��r����N���9�<�cD8Z�����I����3SU�| 84���`GzMUd.���.j�n$En]v�]�QI�$'���8jݰ���vku���U娴�9�oMZ��jr8Y���t�E�*-��(9��B���%����ʫv�R�&���,�3�D���bE�7h�]�T���G;	����ZJ����|xQ�hlY��cRZ��4$EP�2��ܨ���MѸV8�oG�xO��٫o3�y�ԝ�_�2����h(�Wt�C��Q�&�%�T��@$��b�XKW_��|��Tum7'�V�7 �ה 9Һ
�W{���14����6�`����҅���#3��i��D-b:)'A�C��U�èK���֖!�v.���^dXxm��pvrw��q)���e&~m"ᲿL�)Yev[v����'=�M1 V���R����&��M@�y� p"油�ku�=+��(wh��(�"q�������[�G�,p��X5i��!Og���튋�JB\"��t��.���kA����e[��JS	�5I�u_�}�Գ�"!B��[
%n�ʠ�i��B}���d��Le4x�r�B5+�go���Ӥ	2�#QFnb����x����P���ՉM�h�r;v�~W��@Ϥ纳r `��е<�ߘ�`��m^��6tT	�b,-��\JJJ��䉰�$�z%��>Z>h  ��d��~w���6�%Sd��Y(�k�m��x*���[�옧7���`�ڰ�a���کJ�	U�V��@@�`3�=�x$�a���!�X��W���Ո��.9Ȧ��
��,�m��)�4'�� V�u���n���k�0�ۓ�Z��B�]�rpȚ�l�uz�k0�
k���9m�9�/���_JLZyG��N�ǏsX�_Z�t����i<�bR_�*���u�onf!�i/���g����;���x��-�����ʄ���q���9��
p�Hqa�_�'�Ru��(%ۛ>µo�ٗ��U�p������D�%�L��8��.�$=���:6��F>�O��f�ϛ���v(��b
0��4}p�Aa�𰒃P�?��6�b���ij
� �xŹ�Fb�YV����$�L���Ub���(�T��/1鑡U9�7/�¶�CO�K~(t�-�;�: D�L-U��3�l}�A��BwSj�2N�rA��"{`~���b��'��ib@��̓gp)�э>E+�{3e�"f���;Ԛ��ݫ#G�7������5}����ƾ'*�替RIY�Id�pǇ�#}���vz��7���k$X�:�`+���,t !��*�VL�W��	���D5��x,e��<v���:�%[��t�K#����;��*��&l�:S+����)J�_ �y�i$��Dr����5�UE[u)ekry_�5�*�C!�eO4?�ή��D/Ę�6b��:����m=Jg\w��ʡ�c�W�Tw�_����Jæ�.l $!���f�b���M�Re�`OQyf��p=Ț�L�a���%���="����b�q�
�L�]n��t��)c�h�P�j�C�*Y$�;1��Y����I|	臦�&7�~�����e�Q8�Z�d�����J�։.�I�aCP=�AG,�@3K_SR�VZ�\���!��8�Z][4���C;�{��]M�H��b6��l��"s~���*����C��7FV6'n� �_/�*��Ƴ�<W��o#CQ=E7ʕ�P=d��:3^ᆿ2�M&.e���#�&����pq���9`U @�����Wޜ5
6T[��Q�Lz�,罿~q��X�XU��1��['-�º5&��*_,{;П]d-���n/����E��-��T*Dcqͳ:8��gD��6u��^	��֨�Z'#Ղ�R��7�g���B=H���C��;�������m��4�d3Xvf�=cdL�\�v!']rp���7�Eog^��A_gc����E&5xv!1�݂����{�v��ش�y~3�������&��#����0��,iF��eX bx���9�2���,�'�M�h�Ýε��Z��}�v��R_�1<�k 㨅��If�YK=:[%}�,�e�t�_��'9e�ƛ�E��u���M����f���T����_4��SJ�O3]�)m���[�H�|�p0���!!��uT�]�+�����O�Y�"�ۆ� �z��W������� 3�x��PJWl6d?�V�OyK.ߞo�ɽ����ݡ�CV�V�~������� I�A�3������[��gM��bBm�A;k�v���`n�[=���|=9k{�%����y��Z����MC]�%��)i+L��v_,m�%ZA���yvzkcr�%(�v�pl͌e�h����� K����.i���wx=�z��\����sq�:�K��x��H�N�kt��U���>B�WH1%o�X:p��NA�,�j`б�r�eJS��DSF����K�q�%k�-���S��^�ŀ���o�b���o6nh��=��ң��� ��k\�h�C�V�A#\����B��'����m����H��1W?��aD�`.�$}�>n0�9 ���;ļ�B�˔Tl
��*�_��g:	���@�dvX�ߛ%cGK��q���J]�~�4�����W���F�I:��V�B-8pۮ��=�N�_��n}�� y��K.V�� z�M���wU>��g|'ѐ��XeE������h��N--����v:�M˞�P�N���a���ap%�f�[cT��[:�㌰.i{m�̆��w�����8�>�ǽ�1�5;�DVZG�H�ʞ7sm@��|�6a�� �]���hl�(_�c��eO��_�tRR�����A���#ƶ��)���	1F�x�b�9�Ɇ+�a�����V\�lt�<5d�P�8��7G��O
�b`EQ�M)���"�*53��g��j���Yx�8����^�Ku�~��q���B>A�6�Շ)��c��{o
_6s4I�����jK%���@�P4�hɆ�գ	�gzV��Yi�f�,��+�~�(WM�U�G��S��B5źgu��N*����0�s�a�Ч��9خOڒ����z�Լ�����Jq�x����ұ_�:���"-�Pwqa���=�Ң^�lqQ(8Op�9}���aW���Z���,o>6��`�����t�V�D$��G`��sr#ûkv^ ��B�sr�CM6��=?S=��٭'qꭄY;&	�&�1�����|ސ�죺UB+*۷���k��Ɉ()���)��tL%A��Y5	�I��i�)��U��n�?z0��k=#"�u���Ll�F�E���͏��z��i��h�����gS�n�������nU^�����@+�=��k^QN,h��4���AML�4;A,�#8�xD%�u���9J�l���E<�*��[ ��NB�o_��G��6����d�� �n���-������?���C8�p.��3|���ʍI��8)��o��P�k�az��=�o�?S�!�¼�����;�ړ?� �*ϖ�]XAO����V�:	�J��Tzj�nPD)?�͖r����0���3e*g�Y9��~<#󸛼8}����𓮓�ӂ��;vFX�L���F8��:���tE��ZG�c��%#�i������"_�4  >�<6�q��x�����L�T��2�m.E�m��Ts��5��,'��':��Z�N����ۯ��P�~y����ECS�\��������=�N��8����^��I\k�U]j���DsYP�Z��J%�ݴu	�"n�1��e�����`j{�0���h�v�����qD�������O"\�}o�
�T�v�oۃ�&����A�#�(�[�[K�4/�k>m���
�pL�ө�
QYy�#��}19Y�ƖX�6u��Ʋ�����eT'��5�2	ʄ)IU�/j:d(��&�`�q5%�em�/��n�Z���3Mc��b�W$l�}K�!v�.��L4�k[$=��>\a��G��6�<n g(�jMl����	���K�q��z�\�(�؅�w�ŕ��kB���m&]{�`U��loX�BdY�̘m�q/Զ*�����RD*��?`�b�	to�jy+��LoI%�à������yNC���]E*��6w���ۣ3Xn:>���;�sr0ҕd�J=ٻ�^Z�uZ��b�&����T�|%s`O`r��n��{��D�R9PH?P�ł间,t�,z�k��;��HZ,^�{���IK��os��@��l$?�� ��.�_ �p��#�6!�ޥ��$���H�Dr�jz� �#!��S:ʳΊO~��%�{R�&S����O��E��U�Q�ΨSwI���yMte��'G��S�k��aӺKΓ|��@Sb��븠���Ġ�86�?�E7���$�; }1+#��B�C��:6��GL�����}dx�~-dX$cX��'���<a�<!���y�	��Y�t�2��2^��DÊ�]����b�'D�$�c!+���J�i���H�-�*�_L�$Z��׈�8�SX�f�\p�n(���h�P�0��u��kT՛��rQ��Y��7�΅7Cbj��<)QnM�8F2����0�+����2D��r��9�� ~��Pp�7M��$���`"�Q�qM�^������2mZ'�T(=�'��0;NB����$�JRF�&�P��՗r{"rsla����(!KR�[)%�b�APD(�{��ժ�Z�l@p�-Q���%}I_�2������/U���oy��,�<�7�W�QA�#g���{�N���׊	F5�0BI� ]��� >Q6�;Z�kM|�R��K>�(b��5J�>l&m�)�Vr�m���9ڥ�S��L��Bf���SU.��a�J��NÔ�_ߋ8챤9S'��ˊh�x�c��s���i��V���w�Zx�e�zH��On�)HɊj0���,Y��r��@}vӳ�kF7�Z�jCG���Qk㥛F�'��/Z��=��r�
}퇨�w���I/�����1~޹�!�Ђ/C��e�/5. I(�N�^P�/#��6�1���ܵ��X�Ɲ�T�Ht)_I�t�8a�;��י\z�р/�"fP�3�J)wR��%����=jh�`��"y�)ސ�˱w��@�n� ���te
�Z5�C�7���r�P]w
���'�t�b� �G��l1 �e�I�͸,��_���ם���1���z���A������ؿ�EA�c��ƾeLĳh�7~?mc�Ɨ�>�,�U%Q�>�l�̙2�k2�f���}�J��X$\0n�� �c�:B�l�ؗC7�W����I����n{��Y$�qkdUDX��*R4g��[��� �z�w�;@88�dPz#´b.��G�	�*c�jGp�
E��+�T>�wɍTKB��\�����S��g����~�W�s��ೂ���36��giV���7{LP���y�>���h�|Fo�b-�%Y�>B��ݼ��ǆ�z�r��a����7U���[F�T`�^'����N����V�W.������Fb��!i�)��9wڜ*�1����l{J˴!O5�J�ɧ�JTL���Z5��L�����B��Fp��ck�ɫz�y�"Z�Y"���',�] �f�:֞�C�'�sJ8^s�`���#dD�/��-��v�6)�=�i�
�V̮sSK�I�W��`$�һ�~����:��,�x��a�5xP�5ꬽ&���YO��%�Tw^m�V|��H�'���'�=.=��y����/���9b9���3�t̃�rh���7o������׎J�-��`��TS�	:����b�C���3�e,+�HH�zE�nU�^$�Txoݡ�+b���e8V�a�&�y4	B���_��^pPAZKT���k���2��Ò�@��irF�5$C�[�J�2Á]�a�
�fY����9���H9bn�$�T���{��!�
�U��菀@�E���]�8��{֏����0p%�u�Y�U���y����
��w%Z�]���d
��J´�"Tp)+�����㺘�W yF����h/ڎC1ٺ0�����L���D�8}���F��τHr�~�0�R���,�qQ9bX��#H��h�_r�yH�����q�$K�b�)�H�6]��uXdO�>�fæ�;��[���^A�Hr�E�SehM�QP�Yo��t:��|y�k�p��t�<��G��b�x?{��K�X��w"�K� 0���O��hO����u���r�%��գy�vh�{%j��s��P�:� �(1,ִ�!�;`�z�������>:=�
�AY�F�?� ��~(�m�N[��i�(ؒ���S�+��>�ʚC�ԗP��WΡ/��IZv@��գ�2n��̓S4.���F���_�^-
bv����#�O�=��|�k���`b7S�LZ��.zNE��:���)���������?�|(:��	����k��*d�dv�w�� E�Y�A�V�a����Z��tdI��Հ�G�wP�Y��[�_)��93�E�1�����k��>&�n��}��ٽ���������y[�_>�,�LrR7����-� c�b�8S��vGѨFt��(�''�j�1�_F��tW��#�ͮ#��_�.,���f��o:$��_���k��i��H`o�&�����B^5'$+|�K ��Y>�SB-�?N��d����g��������
Q�� g,�AD�Z���<z��r_&�b8~��F����#�g�6j"����%L<'��b�޸� ��ɟ����-wg*���O�#��$�o�ԓ���� hCW��J*�1|	J��؛�������s-B��ø�
FY�A��
����g����86���V�@E���\��@�v�p8��� ��AV�����O!��Ty��-�����@A�CDxd(�5)H��qkcI�؍��}[�]�����AWX\��p�&'��u��n\d�W��xw�i�x�����C侮7%!H�Y,zUkS�ma��Ë�B&�߃5rN�������Gw�<Z�˼��XM3�7�s����P��;�'�Y?�U��H��7C�v��H嶴o��8�	��[î!=.����% �=?�نFg��Ngq=����GB�`t�y�yxɱBs��\���8h2}��0�Ѩ�Q���eu�� @a]�$)\�Bk���W�'{�z���Y;�إ&���z*�!Ĳ�~���X�.��˕�etfn��R�cd*#��<{�&w �3ь�B��"� U3�8�|mf��d9;��%���a'+�E�������8�@yv�V�*��),�b�Uə nP�4�ٿ��E��o�����RY��ꄭ��g�	~fW��x�i����w/��R͕~��'�X��4#�ʍ�H�\i����~U�}I*��3M�E�c�/�p��#]*ȕdˋ���{�H��XM��9�{�@ð
�����[~�FDFּ^q;��[L�v,�Ӽ�ܠ0�H~wM�V+p��1�+�2�)�9H~*�	��`)����2�ūt���2M�@���KO����\�w�!�{����SX�,�u:�d�mfxͼ�{���nʽ[6g�dRsso��l�lx�
�UC0�9���Nz,�hQS߀�ms�m��iVcR���gل��7M��6��5��I�|����߫-b��Ri�"�=�ߡ���DF�3<��N�m`G���f��" �8$�.������È�T���˜Y��baZN
�ՠw�2p��GQ�m:,?��%9���'QM�h��]�.�[e!=֞i�SE�ᄇ-��Xػe���TH0��ܜ���Q����DI"A���*��]ы�0�o���j��r��Lg�54��#a$�*AP��+��`�@��eê�}��i�x�÷!�v/��A�������z�ِ��n��m"F�#�Ɛ	r�^JKob ����Rv|L�<��EG���ӄ��^,o�W/���%ީALg�+WBYK ����֙��,<n �x��`z������V����R��\�+�L�
���	��a����GOm�l�G~�~*�0��.N�w7~;׋>�K�0�r�M67��0�ֈ:�_�"μ��Rg\��6�Ԃp��\X�Z7�1��?�wEq���@`�K��W�=���warUMIYhrD�x�F\���d�^�Wz�л���
>�e�]n��4Z�����%���
�U:̍�-�h��\��ڳ��>��� ����XP�MvX���½�y�!�N���J�,��r���c�AJb�!��E���}����C1]K�7.�X��w��&��m��E����<+6(OOы�Y���0�L�� �f��!�(�<!>�ɹy�w5��i�K��N��2�@	'�M47aր��V�[�����q�hpb����C��l ���U.wG�E#�M&a��9�L\�1�FO��$Z��o�w��+����+w��	�nÔy���|ӈ��RI)6y����'[{0�b�-����XlxV64EB    fa00    2bd0uB�����M!��g79���c+��@��;��%�'���������J!������M--��Ho��<�G����O[�a_S
���j�K����/-H)�D-}¾�ׇ�����:!�>�5ǜ��v�r���ߠGV�,,+�C�>U O��X;��l�>�|��unX�%B�`�g\�Y�x�D�+�������n-D�&�I�=Y{��=�:5.B��v���{���m2N\�l�I��Q���C���Φ#�q�П���z�H�e�w\���p����d�Y?�7��8#lxOO@DKЃ�_��<���̫��S;
l�xwG���"��a�W���7��|��ظ������oJ
��$��7?�Um.���1�*P���.�D���y<>^��d�_�񌍣~Zy�K�=v�CG(=�9W׼���U`��#��~�YX�g,速��b
����7g�� W�;�����xj_�<�p$M�-4Mn���6~�Xu0�1G�׺�?R�M�{n�?�9X&Ŗ�c�vҔ�λ��O�%�a��I-�>n��R-�7@_@;t�6
;�,��5ڝ�!dA�i�s���>�������&/~���I��F��uBIzDZ�
@��d�AHr[�h��!5셌C�ҧ�����"x2���ƒ�[5�C��9�j��s*��L�6�@`�(�v���I+�7�lhX'���y���D�Tu����y�ϲ�g҆���N5vm�G�9��+()H�u�z֎˩�R9	��d�<�B�|�G���bs@ƳAo���e���+k�T�U����݄JH:Ɉ��y�Řl�6|nn�횡�-l�� )_�8FT*a��<��?gŸ��Ň)��y_$_����KP�am��o�&��F�����K��X0Ε�i��Dmz��"�Apx��|G��q3OU4j蕟z=� �A�2��	6�w��{c�lh��DB���g�ݤ~�T5�[�2\�M��ll����<߬��U���V0���I�Z!H�x�k5aY?soK鵀��^�߅e�
�����lp8�G��;.��3߮��_A��)���Gl��qXr�穯���['a(�W��1E;�ewy3�Qj���&�c��_��V��t,���hIfc)�X涙�if'Ϧ��G��Vf�Z
��2����'@�phL[ޫ�^����]�� ~O�	�'����2�??�8�i�8n����?}Z�k��0��{��
��X5���$K"a�#u��Hʸ-�^����X�W����'�p�eot��h(��@ǎ�>��J(�ʟ��HB�B���~DZ:;��Qb���$+�� ���g�j����Iuk�H�Cd�9�_s ��
a�jv��(>T�:�2J:^�7 �1� ���#����㿄PWq%����l���k��冁�:�U��>	%[;nR7�mˬR��'�6$�_բ��_��x���%+,��^e��o,���^�s��n߾�kDx�<�O:�2W�
�f(�l�8]���
Ym^( *bj!�S��ӱ�Ry��s�yEo]��dT�����(�;��(
��}���X�����e��7�8��^J���,8a�'����0:�;ۂ���De?D�eٸ��wk��ɚнh�8�� $�bk����A��^��V/�����kh{��W�-�C#��o�>��uNi��1c����BM�N[l_ÈȘ?g��L����w²���,�74a�4����}�e\1�̀�O��mj��Fc��B0�2���2]%����з7�@�fs��] ���&����="����M��4R���n�O�K��ND��@�ĝ`<9BI��@�V��M�h{~�I��U�c��|�N�!O�f�����g��uQ�j�Ȏ#��Gc�Q�!ys�1��K?#L��Q(o�����:��Z��5ofݨ�T�N�{h^�c���V���3��!�(�r�E%���H�=�����9��Wc�t��H���ᢵ̿g���kJcs�C��e�ѝa��f�4�cY�e���~�yA�Y�AL��]n!���q-���
��l�fə�I#C!o���yᅻ�\��h=`!_`�� �򯃞�O��0B��� �]R������2t���oaP��c�U"jse:��	DRd8�߆fw�+%c���_�m���`e��ܠ{�L��G,�~$CbX����$GT�˾�@�!��5�jlK����i�sD�U.W罳�{�l%�D�@�)�˵��b�߂��q�a�র����1��}�U�P�P5�Q�.j�������%յ���h�����˫qz��%r�|�Ѓ���36�b�FG�ۧ9�l?"�vހ�^�	9�E�����ckWu�͆��Q��]��� �~ �(�3�ѓ��?�}��>�}.�9\d��޸a�zo��� Ɖ��������ɔ�ܚ�Z*�f�n�ls!��Q���U.��������_�$3ҍ�n\z��W�C��_{���RLI��'���xr08�L�;���2�Z ���?넴t��a|���������L7����!<����cJ��;K2�ߦ���~��	��!qhkb��)�� B�P���=X�͚\{ܤ��#ߎf�!.6�к7�^^t3���������'�������S8�$Ж_���%כ�F����v�~��?Mĝ�V�ק}~���i�V�f�7��#2�<�CtP���tU{��eHr�l�;�r�40*���fX��̻��
� `���z�c�3�Ɉ����ޤ 7��*�Ѻk췭��1/�9-����3�0��Ł���K7fYQ_�׼)�~#A=�U��ҥ��!&  �@o�P2;}+Dj������}L�ܚk�$��a�S%>b�C&3�n�Á�F�-Vf���o �;E���Ԫ @�F�,@�reO�%"?�V e>�����'��^ȓ�o�c�-�aM�r����&3^���P�z�<d��nFy!�>� -m���vi��\� �x�!��	SѲ�q�8��G�%t�&�L$4��D�ɲ˵�Q����� t;��^��,|6B�z���Z��+�)C��������P�����J��S\���e���Z��}�<Rl�z8%Q�ɛ�p��Y��1+l�,��U��y�r���Ͼ��$);� ��آ�qk|��`�Ш����,�a�cro���z>�����n�Yr�8�M m�=[�yK-o��I��G�Li;���^oj�BW
�:�^g�Wa���eoU��J�b��s:��n�mʒ���N>��(}�m<о������\)�`u�қ�xu�u� �}�4E�I?{j�M�pLp��%N�0�.�C�T�M_ص��%�����r�7f�3-��=��/��)LrW �*�~ӏX�cx���7�������rT�H_Fm�ͬ;P�m��-��V�^��"Lm�^�H��\�G�E�7�g��F���eЍ�g�x�8�N2���Ty��� D�Pf�R��R��!��LN��;L1������F��Q����+�jJ�k0G�^ 3�,���3 �Md���?�����B��J�����N[|��?���0���!�z`���e����3�U��ư�K|,ߪ7)r�0!���Wz�}�8�
̧Dc\	\4-}��J���&��9_zh���G��kw���P���|�c��u¼�䱕$��*����m.�||�GE�̻��J�?S���xG�~2���q��٦��F"+����y-ݱ{J�����]�+\�-u���(���0�H���j�x4]���A&~(�1��~��B ��y��g$��tل�9�1���ԙ�����G	�g�i��U�r:$ h���20b�hm��d�v7�~X@a�#���JDy^`��6
m�a<E�/ZE�+l�de!���Q��#I��ӯ���}	�j|�4�&��Z�W�eDݭ8����ڱ���D ���&r*5���Iu�L��y�a����
�m�-�_�f��o���^ĶS�N�a�u��Ƴmhqi�'R<���ocy���DߍYH����2�(����0�ԍ�9ƒ��x��čo��n�"��X�8��l;ޗ�! 	���h\ۈH�;��TV�ml��dփ`_y��$ �n�O}R�zS{$x:�����mВ%휙wܤ�����JOWB[ڗ����k�[%�Gf؅C��8���"|\�F1�w^ܻ0E �g,�6Q9��l������=ŽHV=Ƴ��b��&��wuw'����'���&�K������� �QFh״]yE����:O%\Ѩ�����GfȔ����i�*�r�(��H�kw�Da���_1}�艋����li��X�j��3�+I���[Z1��(Ϙ�]��s1CA(��S
���ח����S�被� �+�����퓐HӉtWV���S�ZOP�l#��U� �3�L:&]I~�
$n�&��j/��t�A�S�Ȯ���ٲBX�8%K�_g7OW������'��w��5ΐ��
~��\$�̟L���{�[T�G	�������/����ʄ��8� ���|����e:��Ў�!�m7/��7�m��}~*��%&'�����7V�7؝��O�K����Ed��-E*���4��Zuf����1��z���5K���E ���5�I9����hޟm`�%�jݦ�7%^9�:��d���{���ͳD���ʸm�3C��u��a8����!^������c �����&nrq��Au�;xT�����ބ<qld&*���GP��K�0T�fU�XMR��N��T�=���Є^�t-b�V-H%=��p(x��>c������pv��Be�Zh���O�>���������8�ٰ�/��Ak%ce�J�":����4���wWDd��y`4����-���?�� �ˌI��(^�40�Z�� ǅ渧�YʽJ�M8��vw%H�b�/id�CPȉjy�L�V~�	�}O�!"��	���w��Z�='�H��O$|���
}!�>�7pz��9HK+7W������q�J�u�g=��s����BH�`��a��{gv@�xҀ�GX��ջ{,+bp�jVs�@Ë������.F��*�dnZg���s�������sҵ���=��J�_Z������
H��L��T[V�_�!�)�h����u����eon�J��FԾ��?��.f1�Ϋp�x=|�y���Іw$a⇄�e�n�:��Zzj���ܬ���2���TLb2��l"S$B��$� �&o�u�n�
h��Q�b{�O�DE	����x��P�?U;�����Rαv�,U��[�����7�K�CB��T�i�_k�{ ��I����4*ws�T&d><���y�$�������s:i�3��;�5���Z�k�KWYո�����يA�b�Z�݄��rF%�;�aW�I�ʑ�U�y>���L���'c Wa��\�r�m��Zł;�wF^�@t2yj ���]�*gs����J;'5��f����-栴݅(�6��R�a�ak�	f��U'��+�ި�l�?F�ʴ3Ha�j9m+��sWډ���V%�O@�@h�������[��J�\�Y!�GIG$_�^X�	�-q.�ނd�R��׫�8P<jN�k��M!����W~�y�wE����Ƶ�B����[�᜞Ƣ@���e���c0�_��ޤ�M�l�i�& I?'2r��t��1�������)*1��FI?N����-\L2����`|�89�5�V;�7�c>��l�t��!=2h��)����[a���^T��}�������c�"s�,��TZq	��gitf� f����qy׳Ec����n��K�%�����hoL-�J�_�<O��t��G%pl[��X�]�Z�@E϶#o,kE�ɕ{�mE��p@��w9#j��:����=e���\1�)�Ub�?h�O��ߢ.���
��Zpz�B��m4�p
;��6\�l�x z^�0xr�����ԩ��`����톣����]�cA�D�OP����F*Ϲ�{�&zvE��p�����>l_E�r�j�h�ɍE�ښ�B�S(�ic`��X�Jyqݻ��_Y���Cut��Ck�m�:\�í}��2��-P�Z&W���8����շ[�B
R
t<BVA撣ǖ��LQP���o�+���Y�#��� D�B��B>��b��/U6p/��<\O!/�'ޱ��3��r�$�6o0��Ky�B�a�Х�"|��G�{H.:r��4s�n�)�.3�ѦdO,�!o<4�	��w�M[�+ma�����G�}"l�*զFT{�a�;#�U���J���:l�J����}���Qz��N�\M�dE[2,x����?�4*L��w�8�vquq����Rut�gߏ�����]�f-��5ܠe!����%]����0�E9R ؠ�+��.��]�"���ٳ�&�VOV�ZmM8��ӏ[4B���MPȢp+J0l��
�@
E�Y��Y?�%ԉ������K�`�T�����ߕħ3� ];��vk�Y{Z�x���r��ƿ��{�j!5�tC��n�r��m"�u��E�Ξ�_���y�t���f����Hn�&�m����������t�
L���>[/�+W6�Y��J�V�������x�щ�'�^f���Q���Kâ�r�DVv���L��X"������{�)�=���8�ȫ<�uE�Z�q*�}�Kkm:d:ݓ�b�䀺\��N�SY�L��.T��B�u6�<��f	m>j#3/b��s  ���`�3JH��=~_����fX�����v��:׾LJU=o"?�< T�l����N�~|� �ι�U9(Vp��j�>�/<�gZ´��IQS��e!�����Kf�Hkg]5	��s������7t3m��e[�t4�H�B�3D����(�)���'-��ctm���CDEL-*��d���_�5i*��'9PҤ�?�`?�Ņ��8����\���B9ϲH]�����T=�p �������Mfc��j��C���s��;���p#H��s��'���q���o6�6�S��}� PR�-��[�y��S`b�e��v������0D(��5c;���'pD��ɏ���VmG�@������ev�Zoy�n�l'��M+��ov�?!�s9X9E�ޱo�n��73���'���;:��"�]�2K���)֭/$�^W���^�;�?h����,%g		Y�eo�C�#�-[���֮0-�$��5��kG��I(���^hi����b�}2�)�Y�j�dcH��iì�"�78�SG�&�/c6⶘��� ��m��F�
�U���%.�Jt����G�eEB�ݭ��lXKP���Ҥs]Z�z%����n�Es�&O����E%3�5�RX	���<�	��g<n>����CYO��]M�ّ�_۔Lq�_��?�+;b�����Ҧi$�uQa}��)�y�ޟa��)��/��X�ݽ��ƣ�/�]����T
����^G3+���#��l�k����@gmtY��R�U��8Q��8��9�'q삗+a	�{h��x0�������!��ݪܲ1�x!�o���eĂ�%�����u�����=R<�~�Q|�z�h�saD	Ÿ�#��H�хM��'E�O�I����n,j���W���n�;Z]\:>�ł�U�H�j�li �+�`{��q�#��Y.�p9�p���ICj'W��+2ӇHh��kQ��J ����L���g?�45D���2~�]� �%/&ZǸ�L;S���E��y��K�4���R#��$��8�@[��W�:��,�jkt�}��Z�us$\F����GN揲�/4���g����l	��|��eY��_��P��\�/�<��*��.P�o"�{��&�^��e��b�=S7'�1b��0�.�)���;s�Z���	�-Z��)�y�� ]fi*��A�k�pX ������Y�A�������H���a��ַ&���G��k8n�!�uV��۹vH7u���7����N��pɬ�=
�\�\SG83 �1�}?:�q���[>�����U�&������<:,S
�4�B_^�q?|d-�6�%�a�t:�"��U̩-&�ײ�bIeXnf���){��[��Y_�u�4(л��6�5�)��ٍN�EϹ*f�ϛ ݑ��G�����O��*���o��#�@6��Rʹ�Xɺ����>�T�Ϋq;�Ib��r͖�����ҝ߶	Wpހ�ⷪ��,hS��b���ˈ=d,��8D'���3���x	���Hyu��]�0���{�r�M1k����������M�|��cV�F�_�-�7�-,Ƅ�a��ixww�+2�R�L%��f>K�F�ic[C�"�^(�Z��CC>�ҒrZ��"�P2���4�d>�P�j��?q1z��YUA'�����L��E�s.�������S<��{�̭k����uL}�l�q��~�}�"�M�M����E#���w��M%�~�]�*H�[z��J�6}����i[�I0y��O��`n���gY���/�V�z6IS �L�f�B9�άT���6�/�Q��S��A���MKB8�pFu�I��ð�4>�襇G�շ�ˉ���l� J1y�'r2*������j0k���wR�b�k��EL��z%�byѴ����Q "_��eu�|��wJ
A�
v�{dQQl'�qeuV\恶�~�MhÁ��%)g���Ҹ�+���J�`KT���-��S�WN}.Ň�ʟ��Ś������;�KF�O�2�%Q�^��#ΉԊ����1�]Ri8�)I���DL�P�U/�:6a��֕�JkH$���x>dR'�PB�ϣ�B�n��#�h�+]7^Y���� ����'�O���� �s
Z-/��ό c��%����(!p��+�aE]c�u� �MXH/�O�g�&r�_��UY�47�y����샨ﳖ���!A��ax43i4�=���/ͷ�DB�p��`ߕZ
$ʩ�}j�W��j+���e
��n	-=�=��A|NG9��2������)|��:r��p�F4+@eL������x�exT�4UZ�*�ڤ�2۷����"/�&½���f��uTd
����&G������|���1�V�A 7��.�7@"u�(P`o��(�(nhy�|��'�^*9�@c�`�G vI�ף-sr��\��cN +J!	��D���v��)��Pt��$GPJ��SQ�����B���$/�uP�2|����p�8ǂ�
�F����SN�������u�K�����a?�gY�-�3��:-��&2�i/�6P�M��?��N��Ƽ%$�X��l��������Ɉ�YT�m���R���V�OG向<�+2a:�`t��s��#�1$�D����Հ�()���5����޻5(�̈*q�"w���3�\Y�[2�I�sؘ�yZI��Q���D���m
����C,Gh� l��������:�/	�E����{�{�ݨ?�i� �5 ��!�q�Z �Q6E�<I���#�i�lE�N@��w�?�Z�2��+��y�H��:�#��p��=V�S�:_G(��>�#^3S%�l8���^Z����h3�̼a�Q�r9(j���)}�8�� �m���%�� ��iI��	?����pzg��f����,��`�\�{$�.'}��̕��
K:X�*WL�F}�<]Qr�fӚ3�t��U<*T��hf�k؃HM��9��a���e��?2L�X�J�c��������촡0�m@}P&ôO�l��
Ԇ�zRb�%�������w �c�'�s��8�kw���w����e�1�4�;2G�qV��un��h(�4M�<qS�y�cXL�P� �`j�64�͹{��Y��7�`6"��H�B1�	3P_�85�U^8�ϔ���D5�x̠��/�U�%��ޖ��F^�\/�ʔ�r<*�ձk�W0��M�L�+��q��^)�4��e!��.�j.9A��^�X��/d�\�6"@Y��;M>�[�lX�c؈ZCWئΒ>Sw`Kt!T�=�[�NL�ל�#=w�6-�FN��ڋѮ!��S�Xjs"���v����ݡ��a�����hRU�x�B��ڈ&6�r3�#$���K��ƒ�ָ��z: �Y�P�eo��a����+�	8�� \�U���ӿ2���#g�=ei]j7M�=�`�\n�ݼ���g�aK�j��$���z����=�! ��A�:cq�;�_�AGs�`����y�S�I�W)B�����aa�`�����e�ě���*8�:6��!�:i96�^C�����!AɌ#V�!t�Ԩ�b���*�������SH8߰�({�s?R��ҹm��n�m�b�#=!;v[�r�tz%��{� �(�>�ײ��'��A��Lo�d�B��� xx���H�-}16 �I�R��Y]&uo)���[�B{O�q�����Mص���zNc��!c�O��X��4B�I�l�^��G�l8����#95"A�X}ǜ�?&aw��>�  g�\���| v8>����_!G��3fä[��M���gG{�+��2C;��ǵ���St0�t��U�t�#V��^'�	+*E��� XSY��N5�\g|�pwѷT�B��\z2'��[&7ը}U�������͜�S��F�F·M��O���(������O\���-�I�)���a\�N��/GaM�y��1wEُ���.ɦM_�絚x�ј��}����
���E�{�h]j����P6&y
�� �b��E�V��xm;ϴ���_cl��]o�;�]���%k@�Y�Y��%�p��p!�Gق���{[��ra�7�[�(@w@�ů��J���/�����&GNN����n�*-?gF=LM`͖��M:���"P;~a��0�xr������S�a^�:U����ZB])*2�XlxV64EB    c84c    20f0�)R{q�S�|��Fxhz�ٝ�$13�n�O.	:��&cr8��~��ǧ[�����|�*;��r*l��FJ f|��Ġx���Jݥ��/���T�1K�:j	�#" ����Bh8[2�g�~�Z�)�S���p���_�N7W�����ۯq���#��w0�.�rMc������YX�v��k9��l{��=q|�u	�������غV����Ș��c��ş�������vz���6mJ�t1#��\!�PUVj�q9�B�'8���P��Tf������&S�_ l�!��<.K�����؇�snF��?Y�A�y�R˄�1�Xc�����u�u/�j���8"��ݙ�3�%X�@���[�*!��]-�M��L�Q��L19�T�U�vb$B1��!��u�r�/�x%l��Y���C#�@���qغa	i:�ڣ� A~�8���[��"��/K� ��F����$*{��ea��U;�yI�ߢ��1U�Ӄ�'�$�f�%�Eg"�Ҕ[�V��Q�R��N�Jp3�6�q73����cw�|v^?���$!�a�,p@�$z��Y��oV�<�O4Z%]��Y�>�N�&�$4He~ 	�	_,8��������K���|���DꎄT��0�bT�[���T�99�T��:���t�FHZNH$P�"���[���SO�p��!
�y� �����E|G?��y�����I]y�ƛ|� �zs8���z�,�`Q��Wt�U��쌝A;x�]�����H3�E%��Pn�qG06a��1p��I7���J>:��/u:ۖ�÷*�ӟBW%\8���T�C��d���j�L�RM;�玷H�Ev7����r֋n�6Oe���YO�t���?	��xբ:�ӮW��eܥ�F�K}���t� �Ҝ�$��$��g������LO	v�z�l�Y�f�z��C�8�ѧ�౲�~k�wb���Yd����uv��1/��9U��=��&��ಣ�lB�)�(�
ʤ�����5ݝ���W��ͤE�Z���97R?x�|!v��l���_��hXsrb[��0��kd՛*�R��	_��s�~oK�����]��Ǖ��k��0ʥ)<���,*�k����I�fZ� 3�B�v�ѯ+w7�K�a��\qc�����FL���"��S,����˛�������k��ځjO�N��x���r�w��h���Ka9L��9�j���6���/��۞%<Z��Ép�Q���6H0+=t��$�7�KUC���tQ��$b�Gp"�7���kx����fz������Thv�*)�y��A}��EM�m�d���*�B?OH�A���b!��i����nΪ�nQT��(Äw��)K&�\�'rNؾ�*�я� ��)�.�5v�61U�	R�	P��>���u�։TLu9ɂ
r'�D�.l�B��	x�qDY�6�dǓYۢR�2J��6�0�X����Ͱ�5�\,���p9���;�ƴt�`L�	�
��($�Q�f.�����S1�=3JXK��g9�A�v�3�˪
:�}NRQ�ɺU��m��-�C3����q�� ���+��F�x��U�*���/�AA%O��L�ԬL龜o/�奒E��«��A��}�һ�
������ GWR1�شe�W��"�2�x_c�
�2��w�XL��Qv�X)%ڑ#j��ty#�)��w��c�+�h\+d�N��k{R�����ʶ�mu��5 �D�Ѽ��y��2#�Ua��Ŀk�M�%�3N���DxN\��n� #�!��7��)�N9�&Q����}�/�yR��du��:/�_ d�K�̦%e��7�U�9�D����I�;��qT��l����.G1�膏�O�l�z�H�nD�d"�V���)z�8|M��0����A>9݁�1�&�#e�[��SRV�4���VQp���OT���նH���.ֹ�YP�>�&4� �_P^���6�]E
NЖ���4��B%���Q�D����	�YY�;�B�c[ӆҭ�sx���~��L�P��������Zny��u��2�6�ש�yԆD�����pq���яW2� ,�5~Y�ӱ��]!��X�[{�v���ݰV�A�qC������%�m��!4��S@n�?�ՎO�&��V5r��R��<l朽&~~�����Q���@�z�}��
y&����`���(��D��G'��%�A��/�J��o��J«Eӻ��JCqN�|o6ot�S�w��/�C�/Z��(TM��J6|�D�ǔ[��I��5g<$*��l�}��=�)�=hL"@�Z�;�
Ȝ��N�5;O���6��6�������Y[�_�y/V$NC7U[�y!o�M��I�c��S�+0s@��S4|�5�6``���/����X��h�e��kB���h�w��[�c�}����	vH<�~5�&t�2 ��Իs���.���R�z��w	p�Jt�a���܉��D���7
��sz�����h��ۇ��ǖ�����A_�;(�����S��K��b{[�i��o�T��7��RF4��+�i�x��O�6�g�h����5-Ll6�(�)�-~�v�|љ��	��`�<�YR��xz2�%CB�1��q�l,��	B?��k�I�k�O�������в�����}m���E"rnR�_��*_6�n�/!������d���1���U2��҅Sҟru�q�:���q%=�#�(����+2v�L���P������p+�#�h��Ņ�A�J݄����:�[�"$[w���/���iL?{�=q(�K�q�牳��	,)�@K�;D7+����eBU�q�����\P}�w�)���֛ܩ�2�3	>�ՙ�A�pK�T��涚���cƼGi�<�"k��YA�'��NO�.�L�������M��$K�����^��$C����1��U½���ſ��!��Mݑm���5CI�}�F���a	�x��4�@��D/��	�(}�jWĘ�S��z��+"TCL�,�X�'�I(x��}
k�<4t��ˆ<M�g��e�?6�x�Z��j��v�������O>�]`��k�t4^��݁�l����2�'��1*MV�n{"V��,���@Q�2���ɏ���Y>F�u7�)�sub	�y�ဢ�f>dvR{��P�-����zWƙ��w��/}�(ʖ�	�xd ��)��X�e�B2@	GOy��;D���y�uC\Q��;y�3kِ��@(�ZP�ИV*�X���fJ���*�Tبo��6|z���ר��>|�.�DA�Cɽg�Q�?0�#G �⏨7�F�Jc�����-
�?�5��-Km�/"���Tޙd�8}^��ٯ�*��1]A�~4��,EN�D<���<Z��wJ�nYIz��E�������et�n�&L�T�X6o�(��1��D��4��(�i��jjI�X���$E���m������`�
�Up#^$�a�[�6F�)� �2�X�j�s��9�7���!M�����"3is���E6M���Oed��@��:���ev�E�`nj����)�uaZ�n�д (��cl)N �*_bg���|��8��dm;'���j�'4 eу��4��9��8t���SN�16P��P�%��e�G%�o�����YB���b��Sy���=9��H%��� ����Jd�����7~#;W�z0��\�c�ZêL�k+Ԧ�a8���c��H,���Rm������&V����>��F6�"�t@PI�o|��X=���-�`h�S�}e6C����zkWT/+�8Z���la�63���7���g��+N��R|���ds]�|1��0��g���յ]�?�h}���mo3;�ll�7A��x��
�;C�g�� �J-$c�~|Zl/�$�4W!u؏�V�^��֒�^ә�`���P� -}u!����o\R���`l�*���O��,�? �����cN�����J�	��kz4�����mzޕ������P��Z�
�^��:~�������t�!� �����V�[6�7���Z�����4I�b'K^kp�e�ŀ16��{�ܭ�P;|�Z��ct,W1��w0+ :��4Vs�ML[S�n�c��]���m�(������� �E~J'���M��Mi�Gq��!�!�{�C��8S<L�Ҵx�i-~Y)��/�Ǽ�qE �p�o�OKo/�`Erd���䐞�.�������A�,�a' S`���O��onY�wX
�������~�@�p}���&����78�����8���ɪZ�9���g�MI6
�ӫV��w���ƌ�,�(1�w) ����� a��*G_N���C�����.��ugN)`�x����(�(5���
��宣b�q��H���8ܑ��-�0�����A�@��ω��!-�2����YۏX�6>u#�Ӷ�sO�>Y��]�-e�u��_3���0����q�؃e��>k�f���;c�׾ƫ�&�njQ�Y��Lؔ.�|�Z#�X�E��6�!�J�š��|nŶ�7��FE��J5�  ���!(��&ß�7��� `��z�Z�V��X7a*�ivb���Ba�]]���N(��m8Y�C�^0X=�e�*K|����7m�tE��DT�+Bū쐕���C,O%�N�'[�AV�.˦�xIA���뱫�{D� �j�n�_N�<�1�W��n�oJ��^�zn�ty���bn:<{aS3}�Q�NȖ�]u6�rQ�j/K�g�+[+��~N�b8��"�tsVJ`8�f^���4����s#�{�5���S�)�5�KE�T����D*C'��(�C���S���H�p�* ��	�˪ŉX�C�ƳfyGY�[�OfeԶM�����Co���-⌔s��}D���!���r�b�G��(>����O�oj����ea���qt>��C�*���"'ߤUW��n �P$7�˔<�s��2p���pWÂ��\� �&���>��gearV_�X��>�B�� Z�y�V�o�m�v@�-o� J�����]ʱ1`@cy����Q	���/�ǁL�ȟ�5/l-�NiS8��OF���,C��C��Z���O�X�dOw.��eU_����@�d2���h%Ei�R�E~����Re9f������\F���A�S������b��Ɲ��h��HF�����T>���P���J��0�/{m��D�W�^"��U�w�QZ-xI����V$b�IO��[��[��T�H+�,)��g��w~͘'���v`���=��������c���8i##%J�]E�"�I�m��z �+We{�cȪ��K߉�|�<��0������`�FЍBI�v�E,=� B��#�tQƢ�o�2���?6��Z{8�s �\�NB�@e�%���e����]Tr��\����L�R����1���<(�X/�Ԗ0u��n�u	"�|N�I=�~[�g_�Ŭ;p���y�L�Oz��)g���sh���<�#��R ��%QY~2�ǛWU9�V��a�o�P(����6JG�QU���MV0;ݾPa���3<��p⧷=�5�{_�պ{��i�b�$��1'ܚ�Z)���2����d��3��j���Fm�3�E�v��W��g<*�ũ1��47`����wa�=l����RZ�ƃʹ�Ї�+g���o5���{��� nrJ�l��!�FZ8 ~�0)L�[�Qi���02�V:t1\����T��n>���^�C�١�!Z��R�=���4;�eΙ�Ǯ[//k	ؑ��N �ȴTX-��=8�$���5�eB�'��
v�:����������A��U�2m����Q�;�w���o�9H�u�8"Mm&3Ԫ����ǧ2b՚!k&s]}���m���#�`�F�w�~��H7��i�V4po/�kZv����_��8��J�hH"����K�A��a-	�rp��,����pp��8ׅw�B�������|������J��a���o�@���V���jI��ZBn�۷ b��C����{���5}i���<l���~V��g��Ǭ*&^�u̥.�D���Rs2	ʏ�#Ǘ�I�z���2ק����^c��n�i�^�a7���j��O�x�!9�V��F�&�[���:�$�E8��X��f��Y��+k���IhE��&�a?�'Ni�x�X�_5�4��ԋ=��W2�%���q�Iw��kl�_��Ńȃ��ϑ��8��5\M��WQѶ'V�K֧����,���W����">#AT&!�q�Ko\�e@g�=�'�_��RJ��Dw��4����0��/!K�qޕ��Ӣky���+�B"�� �FP�.m'���'c粒V|����C/N���� (��mʊQ?~�������c�?r�^�"������bd�E�t���-ѷ�5�G|����ٟ�#�Ⱦ��t�\��<H����S>�]�S�{cnڔ�ђ��[G�:6fWٙ���8��T�c��9Y���"~�t����\}��-�r��
JC�k���y�S^k��iޗ�x؏���z��NєK^� �Id��!b�r�!���q�/��;1G������8�XnA�g��R��p��s�~õp��v���'��h�o�>��"º����B��Van�zq�f�~+���� �T�\�4ǿ��L�Ozl�P!E�AI���ؙQY$�A�0-��lҽ�c=&k\q�o3�uQ�	��,�E�N��7�9{Pd'|��z��9�#��ZQEM�9��ݟ�-��?�%ΐ��[?'$�&������1�n�����BW��^L{J0����E\������o4���;�\Î��^{?ZY�)��J��=[���<|�Ҹ�ҧ��N��䠑�4]z��D�Knvç����5p�o�+���
�p�\e=�3��DD-�*0��^�B�Gkҟ��I+_�&��$��Gs�217� �l�m�C�nOwE��95���9�3��>�[�m(���S~����F����@q��[M�X��N�9әN����uf�<�ۗ&:B����"�۞H�=�O3����c�Z���BV�0M��s�׻ t��%���˃��5m�3��KѦ�mp�͸���q�=��F���xcZ���fVp��� �>��h�z��!Q:f
����Z�i����^%c��Ta���Na(E�&������� ��F����2Wl��K'�qæ�m�����5��B��!�*��*�\�5�h��.������iMt�QX\O.6���j[�p�`�+�̨���M��������]��5��ڶ��"�[=�q9�0i���z癛>�s�	m�u`��릋�xFۚ��
���J���ݱ���s��J� ��� E%a�mЋV��=�������tW�{~Fp�[������bP��-�lӛ_9�۔�Q�-�kK��R�����2N�,��կ;e»�4}cz�FB���N��D���	���]��HU���n���0k��g������3ww(ɵr�x�)&�<byJ�v=�G��*���^`���ʦ�� �;�t�{mͺ��>}�6���DQG��MIp����cm�F���qǇ��+����E{�<;�+ �q�ˋ1ї���K�����;kmx�Q�� ��b0�\�HT
���O(E�����RD�Q=�($��3� ��Mm�����)�zC�~۪Gs��ݩU@�̇���ǂ�j�����;e�Ԡ"I�9��w�%��ٶ�8�[/��dO�mG�f�1���{��Bg�����
�EA���_)�}LF�W+I�I)�6j�g���9U���c�'�0�����A?p�+.��m��/A�:�� ��!ր(�@5�&:�)�NnЧ�������W��d���ez{|YmN�ޚ{�Е� ڱ1�ʕj�5��Z�R���&���F]�4X ,J�ad��|;]z��2���5��iU�lrJ��.����a����<H��8���lIu���Vݯ���/�H�7�䲕���5�A��\�Z�'�ؙm@��܂]��<��n����c�۟C�h�X٭�7�߲^Q��6^�؆U~��ک�������$����uZStN_�=�5�"����	<W�1xT���6��F�=���ͺj�v>�uK����	�p1���2tcv˜�0Q(Y��� Y��O(���]>�Q������K?���KA�g�#�sj�b�ɵ��:�Z��8�0�v�88,qĩ�(<�(2jEp�}�cS��