XlxV64EB    fa00    1ec0�Y����
wU4]�I LL��a��Ҟ4~Z�����q�Գ0����o3�Y�'WgX�9NM/�~2-���iQ������6����JG����R�D0*׾� �h�)F�s�6�H�����Ӣ��*F�y��7�D�#��(2�v����K�C�����9�Z���/�aӹ^g�"��B��5���}���L����	(�5�N�="���5���)�E�ys[�{��Ify���c�9�(�fH��=����AN��У�����Z'`iȴ��K�҈�sx!��lZ��X�81M�a����ĀC��2[�lZ�6`M�ى|����^�5��N�^8�����ڨр��(��(��m�@w�J��T�M-x׏�ӀV���<4����~��{}�/;m�r���:&P���L��ŧ�+6�0��p(s�������Uz��u�1��0��&�WK�P����5Ln�\�8Vf#�c��=�u��+:���F؆1�ZL�o	x+C/�±��V�MY��� �p��)�s��:J�6��3�Vy����́��p����^��E�<8֌=٥�Ozр嵕�3)���!��X��d&��Gf �,n�@a�$�y��\b�%Aw5������1�v�pC���s�G�X�*&l�#ڄef;��L+����BfJr8@+�$��id���+�3&=G�Ƨ�:��*-�je"�>�	<�@H��50��IB �ʞ��!i�G�ݟ�P�f�k��UVd�D��/�.<9�۟rq�-Z�c_$a@�ƀbD&W%��!��y�~�o4+yh'�ے|u*���o�xV��tj3؟�|.�	����8�FVTkD����^/k���H��]1�;��KL�U��sb�R(��Z)��
�Q�&m�h�)}��OW/J��8M���pSJ�J��g7I���P��pW���@g�qq���#�v*�V�U���Vf�м���M���%1�_I$��I�|���E�&��F���c�JV�2*/���Fz���ܫe��y�F�p���pL���{~�R=�V�a�|l�"ȟC��������u-3������O�;����^�}T��t��l�����Ćd���>U���ĚV_��S�w̔Fו��������Y��D�-���*�������|US�䇞O�1��p	�O�׃]�A�͠����9�\��f�DX6㽣�m�3CxQ}\^�����%��zm�(��n��)����z�=@���cN�a�vaF��_�"�mcV�u���)E?�vF�n�:od�#�d,�
�Λzt2�2W9-L����܂�A�A��g���I��Qs⛝<�Z�o��*M������z�Uo`I%�D�$��͠���%Ϸַ��jf'��4�I�M�%�Б�c�R���j�m��ձ[͡+s�ѺTIS��~����(�l�5�\*� ����@ZO��)�n8^A��!�P�~,�=X�Mn��S}(� ��6 -��n�;0���MB]�1a+��9�K\\OpX�ޮ\�q���ꝟ�sI�.�ݨD�SX���.��B����W�+=I�- �≑� ���,�DZIl�z��&<���n5q��r䙕C�&���c�}	B'j��]�2��SD+
�O1l�.���ӈ8m��K�;�{�ɟ1f����^7�͗k�r��&�T�s�9�������]�8+���:����(~cr�Gv�(�%�CS6��e R�.��Hۯ�g�U�1;���Ǔ-��Wq6��z�#8��4<����s٨�o\.��`��?T�ʣ���w�gt}�vJ� �%x�|i�	��U+-�p�y�;e�g]4{_�&�swKԞp�v�t%�6U�6�%�eZ2E����M�Zv�1C)��MW����U��;N�BS�Z��n�x�i��4�&:��8�FT�=��\��1s� �(H�G��͋�b�5j�%.\���0�~rq���a���,,��S�u�v��Q��$L��u�LB<�=�?���̍0s ��#��W��Ϝ����"+��7v�l[�N��XO�y�����Yq-��# ��]��h��>�mbyoQ����\�Ok�})�W+ 9�T���t%T�q�m5S^S�+��a˞4�1IKU?q�U�5�(��M��kh[��Z̋{S��,�S�"X�%�2��N[���!�| �т�@�S#�b(.w����*��p��a��-���w8�yGg��WfI�[���k����
I�~�fQR�d�u�:��M��'��>F'��&l��[�� /~�,�x���Z�z���Oo ͼ"��礌
z?�<�oD&���-=q�$���~[Xň[T���G^M4(��P��!P{����T
]JL*�۳E��iI��
��âze�x�Q.3��)�h���&�����r3�V`�Q>�
w�x�ܰZ����wp=U���3,��p%{����b"(=�#F�<�z��W�&�ٝ o��Ǯ=�`�*i��8e�X+H�;�x��=A[w4�	a��l��TE������� !�<k�@P��0�=/�P��+� E{��N%zP��NFj>�K������]��Ț�@*�Ҫ�R�c��A�������у~�u��.�8o�h35�4��h5��E�tN��/Ps.W�,~ny���i��jYљj����Yt�9�	�@�B�p�70�5y�d�F7��X�!R}٠zQ�S/�pK�C�c�:����&v)����q`�Gk��"��*+I�Q�,iNL ���#��U���|1��@G5�'���$%�B,Y;����_�?���(ቕ��!���E%.����ǣJGŇ1B�HШ�<C&	p1N��`x}&�C������щ�
9��$���X��a�ՙ�.���E%/�����\T�x'5
�S����Y߶�������yǨ�6�'P�5�G<KQ�G����Jc��\�i�[�Y���a�s�jhW6p{r��fC��Q�v�GڼiX���h��������t�S�E�O�ho��p��A�ֻ �������n�hʛ��%{^�*�S���?����Z�O��,�м��:511D�jp�eM��bP����ӽZ5n���*�A*�8+pQ;�5V�����5b%D� xU��l�۩ڕD}$�)cɗ;`6���e�|��8�[� �R�0���s#wS�ܰ��$��S��dU��H��B�����0�cCg��͑T�FN�Js�F��o��ڂqK��P`?	��R��*q^v~�K4�Qh�ԥv%`p��M���:U�M���3�!Ij��+�$����#d>�m#ֹT`eYooۣf���3:�K%��]�hCqg�v���Z����Q��ǹ�MW^�Z�
պD0~ݦC�R������`؈��Q�8�6�-�cD��UEZ������4j�8��P}�n��zV��o�����/���3pT��ف�tw�6�50��/��HGB�#��ϗ�����Z;x��̇���aiZxR���-��d��h�1���5)���9�?�]P���s�����G=���c��Ec���p��uU ��~�7��px���'�xt�|�ͬe�]?v��U�f��������%���~<8��mT�^��d�y����ёn����Ʋ)���`r���P
\����Ō��/3j�W[4#�ߚM�q_G��2T��-�����t�x����	=[���2]v ��sxW�Y0���jKy/����ך�{��"�T:�_�(�f�(��=��<�[Q��oG��o/1����H�a20ڪU�9�{�WN�u���޴�{�䟀t�3P���L�\�V���O�C�q����d�{��Kນ�C�4�f�?�`�@_�y��
7����¸V:�C;��YS�!��ݜ	�~�K}���B�I��I�
�~�
����!8q6���-�����/<@N�n�H�:�����f��"��Z��M~��5�UN��1�O�N1z͌�%��Lȟ���7����	;t���=~����{7�Y��!M�h��$��F���Ξ`j�u�nc�f{(�0@�LШ�׻�ܐ����%��eTJ$c��*}�uX {���&7�T=�܉|hM<z���P�ʺ�{}Ɏqd���5�����F\��#e�r>�ƫ��ЖOcM���'�4�8t����Ғ�^���-Di����E'�p�أ������䖌|09x}@r]�B�c:#)����t�Q���mrUU�_I񞃓�������ǅF̥� �D�֨�Sž0��k�E6�qU%�W�1Ҏ�ǃ�,�Z�s�T��7x6	�qW��yb6O���`��FS�s$`����1^�Y$���|��&����������sa�Q�����pF߾w%7�����~]!���q2��ي惣e�1؋�O�cA��S`��};���d�zZ��3lX�g������@䋜�g�%*(�� 9q�~�h����<_��AB�2��D��Yy|���f���5��`!�װ��T;g���rm+�C��|ft�!ܦɁ-��`T�]6�dM�-�c�
G.1p�5u�Β�7�����,"D�P�2���C�G���!<�-�2A��na�_����>#��@�����_��nVٜ�ƽ�t��F�2Pr?#~����a����d�V���+����)��	�2�E=�bBя���@��D�7N�E�m|�9�5��R"��#@;x�9���H�!�J?M����Z<���p�e_v�o)`��y��n�������%���
�Թ-u�<�t�:��O�A6[����z3�RU�x�.Q��m����eF���&l�R�`�w�{�P��Ov���@�%W z)͌^@�n�wܧM����c��,2H�b����1ۂ4��i������Wvq"f��}�"P6J�$�^>`,�L�t�d��9v�Lk��}�q�$U@ԃ��:��bޒ֘?�t+�D9΀p��u�͇�`8�*��9��J��~p�'���c�t���*�g�Gs��)�n���c�����r�7���
m�d�ts����(�>�B�<�|E�ѐ����g�Vʣ;*����3i�dc�L�W>�X�A�����w*�?Յ՘� G]M����)*���k��Ԙ-�׭�?1���{#�˔|Y�����;$ՙ^$�gp��osO�"d�}���\1u|R�sro�2K��;��&A�{���6�8�0�ߵ2=�6h~
��>�om���S2��{Sȇ�|s��������]=�͚q�t*P�Վ�%Y͚��l!g)^��)r�;�4�p\%�y"u��W2Yc2]m�R��HɪzZK���`���MxNC ���*�[zr#�������⶛��c�#
d
�6�n�+�b�K:)dT���������rD��^�KQN��W wy�dfPb����H?)u��n�g�)���琢D�����ooJ�m�T���Up�r�<H�AMS�%� K���&f��{����Jss�\-��O�Uhm��;�����(�{W d���uG���5�Ng~�C6<9�'����-�og;�����:��k<�l���X1b���u�Yn_�(�0��]��&���X�&TH������K_�M̂����_p���CP�����|�q��$���YY��py=:�.5w6_���Zu"y��+(������m.�^��W73�
��f�5��]����}Uܟ�bF��t�Pc��nf�܌4���.��#�_�����/��CL���z�]��n74<�Sa���u��w��5�*aS�bK?m�k��K<cP�]B6�o�8&=��`{ÑQy�o�����)�Y|qGk�<��N6�]va��Dx�\0��9�(�f�v�Xv����!c���*��G�M��ѭ�*b�ˤ�kq�#.��k��iS#�w����U�)�;�$�$�җ�Vʈ-p���_e�C��2Ѣ�r	/��I���6򯂁1I�?{3�K�O�ɣ-�����7&�7f���0A��wWΈ��2��l����ΘE@��L(��VnE�����M�^�)�j'�Om&�mI"�
A��x�̪�j5Ћ@�Y��}��xdq�5�1��%�[�V�Z�!�DLM��N}S�bI�ם*������~�4�q��y}�[�阕�{}��W����/!�W���9S�h�nS��m��R�Bk����d��˙��-�,���~l
��:�D?� �����RG�ɭ�v�v~l\n�����������h˒���,%��#��T'�)�Ϗf�m�w��-�R���$�ul��Wބ2�5k	<S+;g>G�Y����^��7�)��\%�����J�]*8 ��t��3P�A�j:D�U����Ϳl#������R�^+@�3ۀ�%�Z��P�טȣF��?m���G[�1��HV2�����`�b3z�.��o���C�Ҕ�{Y�Q�)V�N�H@��I��Y���t�:Ǘ8RT�c��C����3.BȯH��V43;�l��6�j���)���q&�M���>�h�X��1�܄xXn�s�������ꂊv+[�V��L�O?��P�!�[|�P�@���b��3[d�V���xl���~��8�R��+�YCp�G�}�w�DBD+T�#��n�k��`[��P_�r�����o-�:��B%kmUߔ�M>��aĞ��o���%�~�P���S�X!���ܴʾ����/�����t;���Bv����*�����-G�|���wѾ�a�PJ�D�7���[k�*���Z�ҵE�RA�u�_JP�	;�cw@�����i~y
�VP�/�KF_�ꡔ���R��Avj����R4�s$��y��-�A�>�K����X? �;���[��� �/#[�Լ�ђ}}���j�r���O�I�P�E��iy��
M@��eB�k)�*�E��A4`
H�mϧEjɥ�^��٭I��&��,�,��	����6F��}�sB!�u�꘭?�310��{�����I�@�Si	�SotB��Ss_�p�5-�=�!��Ks�����W��`��6[�ʿ�+p0��.��m{3�m���WQ���=�J�Bbv�n�X�3�s�d6�"P��_��e:G|�:���@��f�	}P�hk;�5�xuЋ�5��`��J�m���8;z|W.z-���+�paXWP�哦��L��XL&�BD���dўa��������䎥e�����s�k�HP�T,<~��$�g3^a���Y�F�D%�a���3a��AD _fB��N�
vCVОm�Tm����b����[�b?5��B%tyz�z?)j;�D2\3�j��b��z��7M-}���06ڨ�`�{��4�3֭(����T�nC5s� t�H��b��a����6bݩ����ᯔ+ݙ
f�U�#ie� �kϞ�C&��<�S��q�i��k�F\�3Jz�Z<#Eo>y'Mޫ�%�D#�t�˕�}�h <e�b���h5J򠳡�����xx�ċd �|_
r�<��v�����6)�ͬ�{j3�o]K��fo��Y{�����6��zU[�$4)B��CM�۶t"7�#���J�]%�8�����E��� �q����j��z��3;d�h�V��z��y�y<&���E����/=E�V�BZ�x��:^h���b31��M.� ��w��}�x?��+�(E�e0�}���W:���~��6�￶XlxV64EB    7bdd     cf0�:��VT�+星���"�K�P�������4a�������W��Hj���_TPt�>!]�B��N�G�֟%1��؈k��ՑG�!�|��%��O�L�M��@�w�Ԁ(�C�S�bw_yTQ�Č��M���}�Յ��:�Qe�l��m�ߛ����=�8_�{r�t�)(�._����mp}Ș�d��qB,�T��o0�pv�/G�A�2�_2�/��.��-��g%��y.:}מ��{���� J�B�«!�v�8�ܚ
���h�u�j�֯��z�R�	5�l��)�یr0��U���b��f��(�!P~�&�$mE��>��˾(�������y����Da��9{t�x��[p�K/�J��Ӵb��A��%I��g[����UYA ���4��vN�eg�����H�d	s�w«NHn��C� ٕ��Z{
���o��Z^����Q�Uk��Q����vm�sY�Bߨ����<�^�!�V�����\���.�A�8���G�]\h��������O�]��?C�x���b]sT�_�f������G+2��Eh��K��A�<��"���R���l���Z��R6Z�_8C���J�-L%K*=��i:�P-�ũT�uh�u�/9�i�M
i����D���˟�P����hp��7��L���� �x{�Kj���R�@"��-"=#�ymo ��*^3��s�-2I�ή'�.w�xO���p�bя�"g��}�հ!d��&l�,뚓6��[0��@��}������l�č�wTxA�">d�a����U��?��?H�cz�{�٭�/*�/ig՚����4| ���Q�9�k�I"�,��
l�ru��ռ���-�V=���j�j�VL�`�x�ҏ�Y�"�O��*-ϔ.6�� z5F�C��1B�G{��sѥAI�<��4���X �߁��HI��8�����Z�[�L'!m�����Ԯu&�"��i���Ƭ����T�e��.WRչ�t#�Cb|�C���W����Ry�I�l+�l-�%1拖rWh`�Yd�ܺ�-�buX�:�Y�JGTp|��B���Lq.��fx*�g��G*�,���~&N��w��򭛄4�B�:�&Iɮ�^J|�6����ρ�"�lۼ��7[6�~-���� YQ�(	Z�y��%s�i�LC{S��!v3�Ӗ��J~ym�+t��LE2��@	X։7�L��p)+�q}Ʉ�qԨUI�(����U�ExM2��=�� 6�,s�Њ@S�` 9�]d�?.(vv6�d��Y���ѥ��� N:w�0��A��m FԎL��Ƨ�4�k�]L��՘�I�mx�����SM�sj(Z�������](y�u�{��92հ��釼憃���X5�{v�Dsԓ10��]D���Ϣ	����A  �S�A���hq�;���X�Y����x����;��`;�@��	�!`�3�}�;8	�|����)k�P�ڸ�Sp�%���FW��!�o�`􅡾n�k�Z�a}��쭐:��X(������"A�[�)�'��$���ya?���;V�g�bվ�^m��ٮ��➳_<��M�.�)�W�J3�<y�W��=kWb~�Ѱk�>�Iu����b�vi�����fۤi����j�>��ly��l7��p:2Õ΄	~��}��"���GR�_����Y����ń�4rGM���| �ҸHy^VV��<�!��'�G
��6YUۡf�ʕ�/������4r,Dg�V�=}��k7�s��qn|4�ŝ����w���3w9�,�w��@�cJ��J�t��\�x��(��?j�w'cj4�]��!�
`�q��(@u�d��wvz��W�E�2��P�0�oTb�����9]g8�f��u>�򪟔�9<�Dm`f��dQ�Cs��=�=4�K�	�m-�ژ�R���k`<	4�;�� ���~P,)���}+4"���9���1c�z�<�9�f�9����NL�UBy~I���=t8"a�����r�D헢�x,`����9'.�,�L�����刃"Dc� eŋAS ô\eweL��ӯyB	gn�dVik���p�?�o���?�6xS]�b�"�U#ƚkc��9���z�^��:߫0�Dc�g�ϗ1��.!�Qy���ٌ�L�)� ��y��"7{�x��ad����=y�*�11`䆲�_b��Yp��;)>�ǼU5�ܠ������< �(�>�>�4�Nӕ.yFp7Q�w�v�BS�m��K���w����g!�"���v�7��vƓ��UŪ7���#��\CY��"=\[	R�0��r�&[n2��О�D:�*�?b���֒�	��Zf�ț1�L��%s�QN��"3;I�ka@�&�s�xV_*Sh�+�4-�u�\Ʀ~$��Bc�7��ʷ�?�tD��ma+�L;ؼ�����Y�D1'�xcYD��Ga��&�
�/M�b��Ҫ��ŕ@J�bO�U ��Ș�H}���ɀ?{%��>1�DP�?�'aE�MҤ�*"Y��͔��ٗ�]�����͂�5��-U|DnU� �a?��G+X�y�1{�	�NA�}��K��t����2z�Pݾ�{:�B�L�����1h�w�w��	�v*�-Ƈa)�}�gӣ=}���`Z`dY��2��s�޸���+�U�@�j[N�n�B��l4e]��#;U�d��F8�Nt�st �-�
��6�V~�R��7I�JEӖk�*V��l�+So�1aP�)D�h"k�t^�g�>������Ȃ���y%�h
c�� �p�[{,�k�g��lC
����OyB��,�����6L�V����Z�nj������,U��"��5NTs���V��wzpΑ��3���ě���
��5I���p�)%�+���[g���c�b����;���ě<�L��O?xD�!��h����-S��	��&�fd����!��^B��B��
Ƶ�=Bo\�ʪen8z����^ob�'�M�d9�b��̶@���G���d����f\R�T���f�9���W\��1��{��t���Ś�.��V�0j.b*z݇E�0Z8�7���񟌅iBn@�b�%�:�f핱m'�i�8����%��y6��/w�����)=������j0���O뤓��f�R�y�>��y�*U��6� o��N�l@C��}���z�>���3���"豠������k��_t(��bA���d�o�ˌp� 	$�f��H��.�/#�EY
�8@��T:��Ph(J*>0��