XlxV64EB    5abc    1270��!S)�rǓ���O�	%'д}$�$\��`�c����'t��W�ʇZ�AV`�G!m�Su���[7�K�/H߽�)�-�4s�"��O�
Q .Y�|�
"��<��͏�&d���b���+�qB���;�OB~�y���-����ޫ��mf�lp�����q�EDqAheZ����7�����}o	��gL�q����P��'\5����ы����.~{��ӂu5��g .�E�������e >���oJK^o�@�䠫q)�͇?:��D�M6���ʔA?����}7����%ղ��y�wC���؀5����-o�Q����?L��EH�+Ƨ:��YT����B�@f1�� M3�^)3˽N���>�V�2�tڒ*䯬�2�=P����\�l�����2R����\p޼Y�~:�[����2�ط���HD����z�O�P�*��a�c ���*��1E���,h��#}���Fl|�9ё��Ǝ
͜�6W���
z�=�\����ʯIik�3L ��CO�Vu-k�Ī-\EB�u�xW:�B�l�u{���0̭I�����М�z���j`�LV=������:�4�((W�2��9L�:���)�O������ _�*1B�*�r��v�.�؇��G�u�8E͓��BY�s�\�����eؒD]�L�o���#����|eê	{`��0P��-�p%�����gv|��,�²=�� ���M��X�*տ�x�����1�m/�g��,�!���D��LK���X����U�c����j0ir*!� ��:�yиsQZ���~U�u�l��GId�ɃQ���/��,�$�2l�T}|�h���}������1�v�խ�������o/�-��0�L�=�6��;�����K#2VeU��9�h׫Ξ���R��Gg@�+��2E�Ҡa�8�((\�Vz&7�����~�\�,F�x��<��K��P(\���1HѨ)��[�'����խ�}�՟��T�oD�!��v*J�P{�sQN �ޗ*�n�����9����V�Z�)����;�����4�{�>�̜^Z��X����uI��ED�c8#�0��mtF��t��V-�d8T�Ce|1��ev�.��E'
!����`�����	Y�dw�h�o��\ L�({&���$�#NA�։�CTX˥�xY����B�o�,*�����F�t�K9(�ż�U6F����$�˥3h����M�����s,�����
VV?�򭪤40	V�Ҕ�)�mͬCW,/�v\�����^}�)E����ʩʘ��v���!&'5�$���O2$��"O����TQj�n�+#�Q�"K��҉��@RpӖu���@��w��B��<��'���a�l�LK3]�/0 |���\8�a�U^�K�b� ˈ�=�ݙԬ����<o!d�T�Z��M}�|��O��U�1<����o��˫m��}�$���Kpֹ>�D�+P���X�=@�Kæ6B"D���7 ���kk�8�c���7wo0{����TM�_/$u�JZ�ik��Y���ʏ�O4������N�^#��77�q]�P�P�"��|�<j�r��"q?�����q �*����Q?!�t��� �e���&`'�̍�D����ۍ��p��>*}��QA��&7�����|X��MI�Գ�&}Q�'�t{�n���\a�XC�k�>Y�<�\��3��E��פ\8Ԭ���A�$��|L(�^>�v�S�ёF�Y5�R#8+"��U�Q  �Ӱ��c�4��71o}��¤�BiCR�>gdf~�=�u����+��=E�J_�����)�W����mh./%(�ԋ���([iۓ��oUS+��>��
y}γ�n�CR��O����C����d�����w�uײ:���U�7��*�('{T�%��(ɨ�S�߭�<
�᮵���{ٶt#�}؍�5��ˌ6��Q��uN�����Y�.����t��T�@��.O����Ҡ��^h�9��qwf~#?�si�	p������>���-x�S_��f����C�A�!��m�>TW}B��z�5�ԋ��^l���%p9Bɨ(���q��نH'<ܟ�ї>�q�l��C���j�K�@j4lgvNel`����B�{օ�(��.x��pq ݵh���L�tʞ׼��z8o�{v5�d�wv/`�ʗg���?�7�L!d���g�=���C'�wm58;���؆+75���&ժy�|��`��M������k�qSN�������M��P�֥�5Y:���ٟ�\��V@�1�w����f���:���M��Y��܏����V��3�Sl�����Xw!�~����[�����oj��6z���3�4C�j���b{��n��Y��i��d,��2K*0�����s'����S{�P��@����;1�y_���U~�V%��p�)�2�0뜳N��s��{���6�	n~E�e��F\A�Q����9��k�ۓT?}��R�{N(�"��4��5+�q2ܻ}�����>�R�GX�/\��Q"����WD��m]���ƭ��GtAqFm��$����P���:Fάv(0����e�9�F���r�r������huxq�^r���cu�D�g���Mć�2��7�UV-x?_���S:���
b��M�b�`zQ����ƪ\#���3���R���`5��yʡʍ?�z�w�=Ҕ��h��bb�P�f����KĽ���&��w�Y����������%I:��ņ`v�o(�ٗS��9e�k�D�c����/B0~���J�᭘R��_��u!�٬������ֹ7��ֲ�rfJ��ݎ�$6s4K�9�#)b��6�b^OD5����[  SjSP��w>�w˴",0-���ov�4gN3]��hܗ�F�*�9c�`2�
)�պ��1�Á�z�}����I?4Ze��Ư�.���]H#���p{9��ϗ����bĕղԸ��X ����LҐ�ب��cnH���� �R�����O��&E��8|R�6�R�/��u�JG�_�Ges��1�m�I#/�P�4m�k��pXK��(�(��mAoN���ΛMI�(-�"���̥�3,(��r�Qa�N�k���j��\�r�$3z&�v��d�\�Ј�n�<��O*+&��K��{sr}6����6�c
��o��_��o�/XQ��gΛ���>qG��d��Zyh�2� lz+v��e
6=��[�r�ti�f=�ܗ Н��<����%ˬ���Z�ކ��%�+r�^���;Ф��Uضؔ� -�������}@�fR�̺�tڰsKB�?��:�����|esl�z��w���4�o����r���7�틊"�V�|�h�?�SB#s����c$�P�a�����y���~��{k��v���v�4NS��<�|i��sIxS��H�A;n�k��p�B���7�Ϲ����t,FQ�N���:��p��7����:��o�Y��HL�)����h��r:'��)�����h����zZ`X�;ʧC\�;5v�f�aG~�I��������!�	�ꆽ[6�*��l�xɞk_��1D��Ȼ
�;�K� ��D��+��c�"���~��ʧ�P&���d���)a�� ����SJ�r���`B3	�q?�fTWE�#���X.KU�Jč�+��D;��Y� b(�T���]sz��s�[S6�z�>:�*Oin� ���)N�Q�H1N���u�Շs4BvĎ 
<��2P���*�r�iDJ�b�ǲΠ�	��2sq��o���T4<�kE��c���]z8�Ei�`Eq���$�I�,&f@�gر�l
5+���A/�,tc(�*�u�W�&�X�R�J)�!H�^�a�����,�=�\�8����R�;�K�NB������^���ú/���
��НԔ�%�� T���u$��"H#mS5EN�G���Kh���y~qU��??H�X��w Ke�$�<=����p}OI0�j�3�Ĉ�G[�j�6��丵8Eq_�=bq��R�f:�[��>:����%W;���y����g�M<��'?6�VT3�J)=Ŵ.*	�9עw+�XM�� ��K����>o-��ջ�p)�OO"��!�j�o�hJ�W��0�%��G��
��Зʮ��
���c��}�쨛{F��߾���.����c���~� �GV>%���J�"q��4e�f�0($x��0�[I`޴۟���>C�Q�j�F�x�P�O"��E&�DI�C) ���2Զ�l�L������ՁR��B��M�H��Py����[�Ri3D��d�F�N���F�O�/U�%�:�N�h�X)@�X<�%B��^3��ɛ�$���?s.H�B�� ��}�me_ ��N�s�6'P�u	��j�5�*ۂ׿���b���:�}=�e��;�\�ԩH�!�9��9���\y�H�TH�'ud��7�p��=��x�޵|�s#|LcJC�JC��G�}-�/�����C�N ���`h�0�`�V�CZ�_1�T}�"E����t'm��q'����hW���ނ�epY����}_��:a�`�:�K�k�(AOU&	��Ts�V򫴄����=���:N��-6�L�M��/)FG�� z�